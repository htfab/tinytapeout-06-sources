magic
tech sky130A
magscale 1 2
timestamp 1707137855
<< viali >>
rect 2145 20553 2179 20587
rect 4905 20553 4939 20587
rect 8125 20553 8159 20587
rect 9505 20553 9539 20587
rect 13553 20553 13587 20587
rect 16129 20553 16163 20587
rect 17049 20553 17083 20587
rect 27169 20553 27203 20587
rect 2789 20485 2823 20519
rect 7481 20485 7515 20519
rect 11713 20485 11747 20519
rect 19441 20485 19475 20519
rect 19809 20485 19843 20519
rect 20453 20485 20487 20519
rect 28089 20485 28123 20519
rect 29990 20485 30024 20519
rect 3433 20417 3467 20451
rect 4721 20417 4755 20451
rect 5825 20417 5859 20451
rect 6009 20417 6043 20451
rect 6561 20417 6595 20451
rect 7573 20417 7607 20451
rect 8309 20417 8343 20451
rect 9689 20417 9723 20451
rect 10425 20417 10459 20451
rect 10885 20417 10919 20451
rect 11989 20417 12023 20451
rect 12173 20417 12207 20451
rect 13737 20417 13771 20451
rect 15209 20417 15243 20451
rect 16313 20417 16347 20451
rect 16865 20417 16899 20451
rect 18705 20417 18739 20451
rect 18889 20417 18923 20451
rect 19901 20417 19935 20451
rect 20361 20417 20395 20451
rect 20545 20417 20579 20451
rect 23305 20417 23339 20451
rect 25605 20417 25639 20451
rect 25697 20417 25731 20451
rect 27353 20417 27387 20451
rect 27813 20417 27847 20451
rect 31585 20417 31619 20451
rect 4261 20349 4295 20383
rect 10149 20349 10183 20383
rect 15301 20349 15335 20383
rect 15485 20349 15519 20383
rect 19533 20349 19567 20383
rect 23213 20349 23247 20383
rect 26065 20349 26099 20383
rect 28641 20349 28675 20383
rect 29745 20349 29779 20383
rect 6745 20281 6779 20315
rect 10333 20281 10367 20315
rect 10425 20281 10459 20315
rect 11069 20281 11103 20315
rect 25881 20281 25915 20315
rect 5917 20213 5951 20247
rect 14841 20213 14875 20247
rect 18797 20213 18831 20247
rect 19625 20213 19659 20247
rect 23673 20213 23707 20247
rect 29193 20213 29227 20247
rect 31125 20213 31159 20247
rect 31677 20213 31711 20247
rect 3433 20009 3467 20043
rect 5365 20009 5399 20043
rect 13553 20009 13587 20043
rect 19993 20009 20027 20043
rect 20177 20009 20211 20043
rect 20637 20009 20671 20043
rect 22109 20009 22143 20043
rect 25881 20009 25915 20043
rect 14565 19941 14599 19975
rect 14933 19941 14967 19975
rect 24593 19941 24627 19975
rect 2145 19873 2179 19907
rect 22937 19873 22971 19907
rect 24869 19873 24903 19907
rect 26801 19873 26835 19907
rect 2605 19805 2639 19839
rect 3249 19805 3283 19839
rect 3985 19805 4019 19839
rect 5917 19805 5951 19839
rect 7113 19805 7147 19839
rect 9137 19805 9171 19839
rect 9393 19805 9427 19839
rect 11069 19805 11103 19839
rect 11713 19805 11747 19839
rect 12265 19805 12299 19839
rect 13737 19805 13771 19839
rect 14749 19805 14783 19839
rect 15025 19805 15059 19839
rect 15485 19805 15519 19839
rect 17325 19805 17359 19839
rect 17581 19805 17615 19839
rect 19533 19805 19567 19839
rect 19625 19805 19659 19839
rect 19983 19805 20017 19839
rect 20821 19805 20855 19839
rect 21097 19805 21131 19839
rect 22017 19805 22051 19839
rect 22201 19805 22235 19839
rect 23029 19805 23063 19839
rect 24961 19805 24995 19839
rect 25697 19805 25731 19839
rect 26709 19805 26743 19839
rect 28089 19805 28123 19839
rect 28549 19805 28583 19839
rect 29745 19805 29779 19839
rect 31585 19805 31619 19839
rect 31861 19805 31895 19839
rect 4230 19737 4264 19771
rect 7358 19737 7392 19771
rect 15752 19737 15786 19771
rect 29193 19737 29227 19771
rect 29990 19737 30024 19771
rect 2789 19669 2823 19703
rect 6101 19669 6135 19703
rect 8493 19669 8527 19703
rect 10517 19669 10551 19703
rect 11161 19669 11195 19703
rect 11805 19669 11839 19703
rect 16865 19669 16899 19703
rect 18705 19669 18739 19703
rect 21005 19669 21039 19703
rect 22661 19669 22695 19703
rect 26341 19669 26375 19703
rect 27905 19669 27939 19703
rect 31125 19669 31159 19703
rect 1777 19465 1811 19499
rect 2421 19465 2455 19499
rect 9137 19465 9171 19499
rect 10517 19465 10551 19499
rect 16037 19465 16071 19499
rect 17049 19465 17083 19499
rect 18613 19465 18647 19499
rect 19901 19465 19935 19499
rect 20453 19465 20487 19499
rect 21373 19465 21407 19499
rect 25421 19465 25455 19499
rect 27169 19465 27203 19499
rect 28365 19465 28399 19499
rect 31677 19465 31711 19499
rect 4414 19397 4448 19431
rect 7849 19397 7883 19431
rect 9289 19397 9323 19431
rect 9505 19397 9539 19431
rect 13829 19397 13863 19431
rect 30542 19397 30576 19431
rect 2237 19329 2271 19363
rect 3065 19329 3099 19363
rect 3249 19329 3283 19363
rect 3341 19329 3375 19363
rect 6837 19329 6871 19363
rect 7021 19329 7055 19363
rect 7665 19329 7699 19363
rect 8309 19329 8343 19363
rect 8493 19329 8527 19363
rect 10425 19329 10459 19363
rect 10885 19329 10919 19363
rect 12081 19329 12115 19363
rect 12357 19329 12391 19363
rect 12817 19329 12851 19363
rect 13185 19329 13219 19363
rect 13553 19329 13587 19363
rect 14657 19329 14691 19363
rect 14924 19329 14958 19363
rect 16865 19329 16899 19363
rect 17877 19329 17911 19363
rect 18061 19329 18095 19363
rect 18797 19329 18831 19363
rect 19441 19329 19475 19363
rect 20361 19329 20395 19363
rect 20637 19329 20671 19363
rect 21281 19329 21315 19363
rect 21465 19329 21499 19363
rect 23213 19329 23247 19363
rect 24225 19329 24259 19363
rect 25237 19329 25271 19363
rect 25421 19329 25455 19363
rect 26341 19329 26375 19363
rect 27537 19329 27571 19363
rect 29478 19329 29512 19363
rect 29745 19329 29779 19363
rect 30297 19329 30331 19363
rect 2881 19261 2915 19295
rect 4169 19261 4203 19295
rect 22201 19261 22235 19295
rect 22293 19261 22327 19295
rect 22385 19261 22419 19295
rect 22477 19261 22511 19295
rect 23121 19261 23155 19295
rect 24317 19261 24351 19295
rect 27445 19261 27479 19295
rect 5549 19193 5583 19227
rect 17969 19193 18003 19227
rect 20821 19193 20855 19227
rect 23581 19193 23615 19227
rect 24593 19193 24627 19227
rect 25881 19193 25915 19227
rect 6929 19125 6963 19159
rect 7481 19125 7515 19159
rect 8677 19125 8711 19159
rect 9321 19125 9355 19159
rect 19533 19125 19567 19159
rect 22017 19125 22051 19159
rect 26065 19125 26099 19159
rect 2973 18921 3007 18955
rect 4169 18921 4203 18955
rect 5549 18921 5583 18955
rect 9229 18921 9263 18955
rect 18705 18921 18739 18955
rect 18797 18921 18831 18955
rect 21189 18921 21223 18955
rect 26525 18921 26559 18955
rect 27353 18921 27387 18955
rect 28089 18921 28123 18955
rect 29009 18921 29043 18955
rect 2789 18853 2823 18887
rect 4261 18853 4295 18887
rect 11713 18853 11747 18887
rect 17233 18853 17267 18887
rect 19717 18853 19751 18887
rect 22385 18853 22419 18887
rect 23581 18853 23615 18887
rect 26985 18853 27019 18887
rect 4629 18785 4663 18819
rect 12449 18785 12483 18819
rect 14841 18785 14875 18819
rect 15209 18785 15243 18819
rect 18889 18785 18923 18819
rect 19901 18785 19935 18819
rect 21925 18785 21959 18819
rect 26065 18785 26099 18819
rect 2145 18717 2179 18751
rect 2329 18717 2363 18751
rect 3341 18717 3375 18751
rect 5641 18717 5675 18751
rect 6285 18717 6319 18751
rect 8217 18717 8251 18751
rect 9137 18717 9171 18751
rect 9505 18717 9539 18751
rect 9597 18717 9631 18751
rect 10977 18717 11011 18751
rect 11621 18717 11655 18751
rect 12173 18717 12207 18751
rect 13369 18717 13403 18751
rect 13461 18717 13495 18751
rect 13553 18717 13587 18751
rect 15025 18717 15059 18751
rect 15669 18717 15703 18751
rect 15853 18717 15887 18751
rect 16681 18717 16715 18751
rect 17141 18717 17175 18751
rect 17325 18717 17359 18751
rect 18613 18717 18647 18751
rect 20545 18717 20579 18751
rect 20638 18717 20672 18751
rect 20821 18717 20855 18751
rect 21051 18717 21085 18751
rect 22017 18717 22051 18751
rect 23305 18717 23339 18751
rect 24593 18717 24627 18751
rect 24777 18717 24811 18751
rect 25421 18717 25455 18751
rect 26157 18717 26191 18751
rect 27445 18717 27479 18751
rect 28273 18717 28307 18751
rect 28825 18717 28859 18751
rect 31217 18717 31251 18751
rect 31677 18717 31711 18751
rect 6193 18649 6227 18683
rect 7972 18649 8006 18683
rect 10793 18649 10827 18683
rect 11161 18649 11195 18683
rect 19441 18649 19475 18683
rect 20913 18649 20947 18683
rect 23581 18649 23615 18683
rect 24685 18649 24719 18683
rect 30950 18649 30984 18683
rect 2237 18581 2271 18615
rect 2973 18581 3007 18615
rect 6837 18581 6871 18615
rect 9781 18581 9815 18615
rect 13185 18581 13219 18615
rect 16037 18581 16071 18615
rect 16497 18581 16531 18615
rect 23397 18581 23431 18615
rect 25329 18581 25363 18615
rect 29837 18581 29871 18615
rect 31769 18581 31803 18615
rect 2605 18377 2639 18411
rect 3709 18377 3743 18411
rect 7179 18377 7213 18411
rect 8033 18377 8067 18411
rect 9045 18377 9079 18411
rect 10793 18377 10827 18411
rect 12725 18377 12759 18411
rect 15117 18377 15151 18411
rect 20637 18377 20671 18411
rect 22109 18377 22143 18411
rect 22753 18377 22787 18411
rect 24593 18377 24627 18411
rect 26433 18377 26467 18411
rect 7389 18309 7423 18343
rect 8217 18309 8251 18343
rect 8861 18309 8895 18343
rect 9965 18309 9999 18343
rect 29368 18309 29402 18343
rect 2145 18241 2179 18275
rect 2329 18241 2363 18275
rect 3065 18241 3099 18275
rect 3525 18241 3559 18275
rect 4436 18241 4470 18275
rect 8125 18241 8159 18275
rect 9137 18241 9171 18275
rect 11069 18241 11103 18275
rect 11161 18241 11195 18275
rect 12265 18241 12299 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 13461 18241 13495 18275
rect 14289 18241 14323 18275
rect 14841 18241 14875 18275
rect 15117 18241 15151 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 16129 18241 16163 18275
rect 20177 18241 20211 18275
rect 22017 18241 22051 18275
rect 22201 18241 22235 18275
rect 22661 18241 22695 18275
rect 22845 18241 22879 18275
rect 24041 18241 24075 18275
rect 24501 18241 24535 18275
rect 24685 18241 24719 18275
rect 25145 18241 25179 18275
rect 26065 18241 26099 18275
rect 27445 18241 27479 18275
rect 28089 18241 28123 18275
rect 2237 18173 2271 18207
rect 2421 18173 2455 18207
rect 3341 18173 3375 18207
rect 4169 18173 4203 18207
rect 19257 18173 19291 18207
rect 25973 18173 26007 18207
rect 29101 18173 29135 18207
rect 30941 18173 30975 18207
rect 7021 18105 7055 18139
rect 8401 18105 8435 18139
rect 8861 18105 8895 18139
rect 13645 18105 13679 18139
rect 15025 18105 15059 18139
rect 19533 18105 19567 18139
rect 30481 18105 30515 18139
rect 3157 18037 3191 18071
rect 5549 18037 5583 18071
rect 7205 18037 7239 18071
rect 7849 18037 7883 18071
rect 10057 18037 10091 18071
rect 11161 18037 11195 18071
rect 13461 18037 13495 18071
rect 14197 18037 14231 18071
rect 15577 18037 15611 18071
rect 16037 18037 16071 18071
rect 19717 18037 19751 18071
rect 20269 18037 20303 18071
rect 23857 18037 23891 18071
rect 25329 18037 25363 18071
rect 27261 18037 27295 18071
rect 28641 18037 28675 18071
rect 31585 18037 31619 18071
rect 2329 17833 2363 17867
rect 2973 17833 3007 17867
rect 3341 17833 3375 17867
rect 4445 17833 4479 17867
rect 11437 17833 11471 17867
rect 12173 17833 12207 17867
rect 19993 17833 20027 17867
rect 23489 17833 23523 17867
rect 2513 17765 2547 17799
rect 4077 17765 4111 17799
rect 7021 17765 7055 17799
rect 10609 17765 10643 17799
rect 11713 17765 11747 17799
rect 15025 17765 15059 17799
rect 14749 17697 14783 17731
rect 16221 17697 16255 17731
rect 19533 17697 19567 17731
rect 19625 17697 19659 17731
rect 26525 17697 26559 17731
rect 3249 17629 3283 17663
rect 3341 17629 3375 17663
rect 3985 17629 4019 17663
rect 4201 17629 4235 17663
rect 5549 17629 5583 17663
rect 6929 17629 6963 17663
rect 7113 17629 7147 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9321 17629 9355 17663
rect 9781 17629 9815 17663
rect 9965 17629 9999 17663
rect 10609 17629 10643 17663
rect 10793 17629 10827 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 12357 17623 12391 17657
rect 12725 17629 12759 17663
rect 12817 17629 12851 17663
rect 13553 17629 13587 17663
rect 14933 17629 14967 17663
rect 15117 17629 15151 17663
rect 15209 17629 15243 17663
rect 15945 17629 15979 17663
rect 16129 17629 16163 17663
rect 16313 17629 16347 17663
rect 16497 17629 16531 17663
rect 17233 17629 17267 17663
rect 17325 17629 17359 17663
rect 17509 17629 17543 17663
rect 17601 17629 17635 17663
rect 18426 17629 18460 17663
rect 18797 17629 18831 17663
rect 18889 17629 18923 17663
rect 19717 17629 19751 17663
rect 19809 17629 19843 17663
rect 23305 17629 23339 17663
rect 23397 17629 23431 17663
rect 26065 17629 26099 17663
rect 28641 17629 28675 17663
rect 31309 17629 31343 17663
rect 31769 17629 31803 17663
rect 2145 17561 2179 17595
rect 6101 17561 6135 17595
rect 7573 17561 7607 17595
rect 7757 17561 7791 17595
rect 8493 17561 8527 17595
rect 12449 17561 12483 17595
rect 12541 17561 12575 17595
rect 13369 17561 13403 17595
rect 13737 17561 13771 17595
rect 15761 17561 15795 17595
rect 23581 17561 23615 17595
rect 24961 17561 24995 17595
rect 26770 17561 26804 17595
rect 31064 17561 31098 17595
rect 2345 17493 2379 17527
rect 5365 17493 5399 17527
rect 6377 17493 6411 17527
rect 9137 17493 9171 17527
rect 9781 17493 9815 17527
rect 17785 17493 17819 17527
rect 18245 17493 18279 17527
rect 18429 17493 18463 17527
rect 23121 17493 23155 17527
rect 24685 17493 24719 17527
rect 25881 17493 25915 17527
rect 27905 17493 27939 17527
rect 28825 17493 28859 17527
rect 29929 17493 29963 17527
rect 31953 17493 31987 17527
rect 3341 17289 3375 17323
rect 5457 17289 5491 17323
rect 6929 17289 6963 17323
rect 9505 17289 9539 17323
rect 12725 17289 12759 17323
rect 12909 17289 12943 17323
rect 13921 17289 13955 17323
rect 15761 17289 15795 17323
rect 18337 17289 18371 17323
rect 18705 17289 18739 17323
rect 19809 17289 19843 17323
rect 20269 17289 20303 17323
rect 25053 17289 25087 17323
rect 26617 17289 26651 17323
rect 2973 17221 3007 17255
rect 6837 17221 6871 17255
rect 8392 17221 8426 17255
rect 10425 17221 10459 17255
rect 12357 17221 12391 17255
rect 12633 17221 12667 17255
rect 23388 17221 23422 17255
rect 29561 17221 29595 17255
rect 30542 17221 30576 17255
rect 3203 17187 3237 17221
rect 2329 17153 2363 17187
rect 4077 17153 4111 17187
rect 4344 17153 4378 17187
rect 10241 17153 10275 17187
rect 10885 17153 10919 17187
rect 11069 17153 11103 17187
rect 11713 17153 11747 17187
rect 12541 17153 12575 17187
rect 13369 17153 13403 17187
rect 13461 17153 13495 17187
rect 13645 17153 13679 17187
rect 13745 17153 13779 17187
rect 14749 17153 14783 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 16313 17153 16347 17187
rect 17693 17153 17727 17187
rect 17877 17153 17911 17187
rect 18521 17153 18555 17187
rect 18797 17153 18831 17187
rect 19441 17153 19475 17187
rect 20729 17153 20763 17187
rect 21281 17153 21315 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 25237 17153 25271 17187
rect 25513 17153 25547 17187
rect 26065 17153 26099 17187
rect 26249 17153 26283 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 28558 17153 28592 17187
rect 29837 17153 29871 17187
rect 2513 17085 2547 17119
rect 7113 17085 7147 17119
rect 7205 17085 7239 17119
rect 8125 17085 8159 17119
rect 11805 17085 11839 17119
rect 15025 17085 15059 17119
rect 19349 17085 19383 17119
rect 23121 17085 23155 17119
rect 25421 17085 25455 17119
rect 28825 17085 28859 17119
rect 30297 17085 30331 17119
rect 15301 17017 15335 17051
rect 21373 17017 21407 17051
rect 24501 17017 24535 17051
rect 2145 16949 2179 16983
rect 3157 16949 3191 16983
rect 7021 16949 7055 16983
rect 10057 16949 10091 16983
rect 10977 16949 11011 16983
rect 15117 16949 15151 16983
rect 17785 16949 17819 16983
rect 20453 16949 20487 16983
rect 22017 16949 22051 16983
rect 25237 16949 25271 16983
rect 27445 16949 27479 16983
rect 31677 16949 31711 16983
rect 8401 16745 8435 16779
rect 12541 16745 12575 16779
rect 14565 16745 14599 16779
rect 15025 16745 15059 16779
rect 15945 16745 15979 16779
rect 21373 16745 21407 16779
rect 24777 16745 24811 16779
rect 27353 16745 27387 16779
rect 31125 16745 31159 16779
rect 2329 16677 2363 16711
rect 7297 16677 7331 16711
rect 8585 16677 8619 16711
rect 12817 16677 12851 16711
rect 16405 16677 16439 16711
rect 28273 16677 28307 16711
rect 2973 16609 3007 16643
rect 3065 16609 3099 16643
rect 3157 16609 3191 16643
rect 3249 16609 3283 16643
rect 3985 16609 4019 16643
rect 5917 16609 5951 16643
rect 9597 16609 9631 16643
rect 9689 16609 9723 16643
rect 9781 16609 9815 16643
rect 10425 16609 10459 16643
rect 10885 16609 10919 16643
rect 12909 16609 12943 16643
rect 14657 16609 14691 16643
rect 15485 16609 15519 16643
rect 20177 16609 20211 16643
rect 22017 16609 22051 16643
rect 29745 16609 29779 16643
rect 2053 16541 2087 16575
rect 2145 16541 2179 16575
rect 9505 16541 9539 16575
rect 10609 16541 10643 16575
rect 10793 16541 10827 16575
rect 11897 16541 11931 16575
rect 12081 16541 12115 16575
rect 12725 16541 12759 16575
rect 13001 16541 13035 16575
rect 13185 16541 13219 16575
rect 14841 16541 14875 16575
rect 15577 16541 15611 16575
rect 15761 16541 15795 16575
rect 16405 16541 16439 16575
rect 16497 16541 16531 16575
rect 17509 16541 17543 16575
rect 17693 16541 17727 16575
rect 19993 16541 20027 16575
rect 22273 16541 22307 16575
rect 23857 16541 23891 16575
rect 24041 16541 24075 16575
rect 24777 16541 24811 16575
rect 24869 16541 24903 16575
rect 28457 16541 28491 16575
rect 28825 16541 28859 16575
rect 30001 16541 30035 16575
rect 31861 16541 31895 16575
rect 2329 16473 2363 16507
rect 4252 16473 4286 16507
rect 6162 16473 6196 16507
rect 8217 16473 8251 16507
rect 14565 16473 14599 16507
rect 16681 16473 16715 16507
rect 19809 16473 19843 16507
rect 21005 16473 21039 16507
rect 21189 16473 21223 16507
rect 25053 16473 25087 16507
rect 26065 16473 26099 16507
rect 28549 16473 28583 16507
rect 28641 16473 28675 16507
rect 2789 16405 2823 16439
rect 5365 16405 5399 16439
rect 8427 16405 8461 16439
rect 9965 16405 9999 16439
rect 12081 16405 12115 16439
rect 17509 16405 17543 16439
rect 19625 16405 19659 16439
rect 19901 16405 19935 16439
rect 23397 16405 23431 16439
rect 23949 16405 23983 16439
rect 24593 16405 24627 16439
rect 31677 16405 31711 16439
rect 1593 16201 1627 16235
rect 2881 16201 2915 16235
rect 3065 16201 3099 16235
rect 4261 16201 4295 16235
rect 5089 16201 5123 16235
rect 10241 16201 10275 16235
rect 15209 16201 15243 16235
rect 16865 16201 16899 16235
rect 18639 16201 18673 16235
rect 19717 16201 19751 16235
rect 20085 16201 20119 16235
rect 23029 16201 23063 16235
rect 25421 16201 25455 16235
rect 27721 16201 27755 16235
rect 29745 16201 29779 16235
rect 31769 16201 31803 16235
rect 3525 16133 3559 16167
rect 5273 16133 5307 16167
rect 5733 16133 5767 16167
rect 9597 16133 9631 16167
rect 14657 16133 14691 16167
rect 15577 16133 15611 16167
rect 16221 16133 16255 16167
rect 18429 16133 18463 16167
rect 19901 16133 19935 16167
rect 20821 16133 20855 16167
rect 22845 16133 22879 16167
rect 23857 16133 23891 16167
rect 2513 16065 2547 16099
rect 3709 16065 3743 16099
rect 3801 16065 3835 16099
rect 4445 16065 4479 16099
rect 4997 16065 5031 16099
rect 6009 16065 6043 16099
rect 6653 16065 6687 16099
rect 6745 16065 6779 16099
rect 11713 16065 11747 16099
rect 11989 16065 12023 16099
rect 13001 16065 13035 16099
rect 15393 16065 15427 16099
rect 15669 16065 15703 16099
rect 16313 16065 16347 16099
rect 17049 16065 17083 16099
rect 17233 16065 17267 16099
rect 19993 16065 20027 16099
rect 20729 16065 20763 16099
rect 20913 16065 20947 16099
rect 25237 16065 25271 16099
rect 26065 16065 26099 16099
rect 26341 16065 26375 16099
rect 27353 16065 27387 16099
rect 28273 16065 28307 16099
rect 29009 16065 29043 16099
rect 29193 16065 29227 16099
rect 30869 16065 30903 16099
rect 31585 16065 31619 16099
rect 3525 15997 3559 16031
rect 5733 15997 5767 16031
rect 6929 15997 6963 16031
rect 11897 15997 11931 16031
rect 17325 15997 17359 16031
rect 24961 15997 24995 16031
rect 25881 15997 25915 16031
rect 27445 15997 27479 16031
rect 31125 15997 31159 16031
rect 5273 15929 5307 15963
rect 5917 15929 5951 15963
rect 10057 15929 10091 15963
rect 10609 15929 10643 15963
rect 20269 15929 20303 15963
rect 22477 15929 22511 15963
rect 25053 15929 25087 15963
rect 29101 15929 29135 15963
rect 2881 15861 2915 15895
rect 8309 15861 8343 15895
rect 10241 15861 10275 15895
rect 11805 15861 11839 15895
rect 12173 15861 12207 15895
rect 18613 15861 18647 15895
rect 18797 15861 18831 15895
rect 22845 15861 22879 15895
rect 23581 15861 23615 15895
rect 28457 15861 28491 15895
rect 6101 15657 6135 15691
rect 8033 15657 8067 15691
rect 9321 15657 9355 15691
rect 11345 15657 11379 15691
rect 15117 15657 15151 15691
rect 15945 15657 15979 15691
rect 17049 15657 17083 15691
rect 17785 15657 17819 15691
rect 18705 15657 18739 15691
rect 21097 15657 21131 15691
rect 21189 15657 21223 15691
rect 21833 15657 21867 15691
rect 23213 15657 23247 15691
rect 25053 15657 25087 15691
rect 28641 15657 28675 15691
rect 30481 15657 30515 15691
rect 31033 15657 31067 15691
rect 13185 15589 13219 15623
rect 14381 15589 14415 15623
rect 18889 15589 18923 15623
rect 28825 15589 28859 15623
rect 2697 15521 2731 15555
rect 7481 15521 7515 15555
rect 12541 15521 12575 15555
rect 13737 15521 13771 15555
rect 21281 15521 21315 15555
rect 23397 15521 23431 15555
rect 23674 15521 23708 15555
rect 28273 15521 28307 15555
rect 2605 15453 2639 15487
rect 3433 15453 3467 15487
rect 8217 15453 8251 15487
rect 10701 15453 10735 15487
rect 12173 15453 12207 15487
rect 12357 15453 12391 15487
rect 12725 15453 12759 15487
rect 13461 15453 13495 15487
rect 14841 15453 14875 15487
rect 15577 15453 15611 15487
rect 15761 15453 15795 15487
rect 16865 15453 16899 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 19717 15453 19751 15487
rect 20545 15453 20579 15487
rect 21005 15453 21039 15487
rect 22017 15453 22051 15487
rect 22201 15453 22235 15487
rect 23489 15453 23523 15487
rect 23581 15453 23615 15487
rect 25237 15453 25271 15487
rect 25329 15453 25363 15487
rect 25421 15453 25455 15487
rect 25513 15453 25547 15487
rect 26065 15453 26099 15487
rect 29745 15453 29779 15487
rect 29929 15453 29963 15487
rect 30389 15463 30423 15497
rect 30573 15453 30607 15487
rect 31217 15453 31251 15487
rect 1777 15385 1811 15419
rect 7236 15385 7270 15419
rect 10434 15385 10468 15419
rect 11313 15385 11347 15419
rect 11529 15385 11563 15419
rect 13369 15385 13403 15419
rect 14381 15385 14415 15419
rect 14933 15385 14967 15419
rect 17969 15385 18003 15419
rect 18521 15385 18555 15419
rect 21741 15385 21775 15419
rect 28641 15385 28675 15419
rect 29837 15385 29871 15419
rect 2237 15317 2271 15351
rect 3341 15317 3375 15351
rect 11161 15317 11195 15351
rect 13553 15317 13587 15351
rect 17601 15317 17635 15351
rect 17769 15317 17803 15351
rect 18731 15317 18765 15351
rect 19901 15317 19935 15351
rect 20361 15317 20395 15351
rect 22385 15317 22419 15351
rect 27537 15317 27571 15351
rect 8217 15113 8251 15147
rect 16129 15113 16163 15147
rect 17049 15113 17083 15147
rect 18521 15113 18555 15147
rect 22293 15113 22327 15147
rect 24685 15113 24719 15147
rect 27169 15113 27203 15147
rect 28365 15113 28399 15147
rect 29469 15113 29503 15147
rect 8953 15045 8987 15079
rect 9413 15045 9447 15079
rect 10517 15045 10551 15079
rect 16313 15045 16347 15079
rect 17601 15045 17635 15079
rect 19533 15045 19567 15079
rect 20605 15045 20639 15079
rect 20821 15045 20855 15079
rect 24133 15045 24167 15079
rect 27321 15045 27355 15079
rect 27537 15045 27571 15079
rect 27997 15045 28031 15079
rect 28213 15045 28247 15079
rect 2513 14977 2547 15011
rect 3525 14977 3559 15011
rect 6929 14977 6963 15011
rect 8033 14977 8067 15011
rect 8677 14977 8711 15011
rect 8769 14977 8803 15011
rect 9689 14977 9723 15011
rect 13185 14977 13219 15011
rect 13645 14977 13679 15011
rect 13921 14977 13955 15011
rect 14473 14977 14507 15011
rect 15117 14977 15151 15011
rect 15301 14977 15335 15011
rect 15393 14977 15427 15011
rect 16037 14977 16071 15011
rect 16865 14977 16899 15011
rect 16957 14977 16991 15011
rect 17141 14977 17175 15011
rect 17785 14977 17819 15011
rect 17969 14977 18003 15011
rect 18061 14977 18095 15011
rect 19901 14977 19935 15011
rect 19993 14977 20027 15011
rect 22385 14977 22419 15011
rect 22477 14977 22511 15011
rect 22845 14977 22879 15011
rect 23213 14977 23247 15011
rect 23857 14977 23891 15011
rect 23949 14977 23983 15011
rect 24961 14977 24995 15011
rect 25789 14977 25823 15011
rect 26065 14977 26099 15011
rect 29377 14977 29411 15011
rect 31410 14977 31444 15011
rect 31677 14977 31711 15011
rect 2605 14909 2639 14943
rect 3617 14909 3651 14943
rect 7205 14909 7239 14943
rect 9413 14909 9447 14943
rect 14105 14909 14139 14943
rect 18705 14909 18739 14943
rect 18797 14909 18831 14943
rect 18889 14909 18923 14943
rect 18981 14909 19015 14943
rect 19625 14909 19659 14943
rect 19717 14909 19751 14943
rect 25697 14909 25731 14943
rect 26157 14909 26191 14943
rect 29745 14909 29779 14943
rect 2881 14841 2915 14875
rect 7021 14841 7055 14875
rect 10149 14841 10183 14875
rect 20453 14841 20487 14875
rect 30297 14841 30331 14875
rect 3801 14773 3835 14807
rect 7113 14773 7147 14807
rect 8953 14773 8987 14807
rect 9597 14773 9631 14807
rect 10517 14773 10551 14807
rect 10701 14773 10735 14807
rect 15393 14773 15427 14807
rect 15577 14773 15611 14807
rect 16313 14773 16347 14807
rect 20637 14773 20671 14807
rect 23673 14773 23707 14807
rect 23857 14773 23891 14807
rect 25513 14773 25547 14807
rect 27353 14773 27387 14807
rect 28181 14773 28215 14807
rect 29653 14773 29687 14807
rect 29837 14773 29871 14807
rect 4169 14569 4203 14603
rect 8401 14569 8435 14603
rect 9965 14569 9999 14603
rect 10517 14569 10551 14603
rect 12725 14569 12759 14603
rect 13277 14569 13311 14603
rect 13553 14569 13587 14603
rect 21189 14569 21223 14603
rect 24777 14569 24811 14603
rect 25145 14569 25179 14603
rect 26893 14569 26927 14603
rect 6469 14501 6503 14535
rect 2697 14433 2731 14467
rect 7849 14433 7883 14467
rect 11897 14433 11931 14467
rect 14289 14433 14323 14467
rect 16865 14433 16899 14467
rect 22201 14433 22235 14467
rect 26801 14433 26835 14467
rect 26985 14433 27019 14467
rect 29745 14433 29779 14467
rect 2605 14365 2639 14399
rect 6653 14365 6687 14399
rect 6745 14365 6779 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 8585 14365 8619 14399
rect 9505 14365 9539 14399
rect 9781 14365 9815 14399
rect 12449 14365 12483 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 14545 14365 14579 14399
rect 16129 14365 16163 14399
rect 17121 14365 17155 14399
rect 19809 14365 19843 14399
rect 20076 14365 20110 14399
rect 22477 14365 22511 14399
rect 22661 14365 22695 14399
rect 23213 14365 23247 14399
rect 23673 14365 23707 14399
rect 24777 14365 24811 14399
rect 24961 14365 24995 14399
rect 25605 14365 25639 14399
rect 25698 14365 25732 14399
rect 25881 14365 25915 14399
rect 26089 14365 26123 14399
rect 26709 14365 26743 14399
rect 28273 14365 28307 14399
rect 28917 14365 28951 14399
rect 30001 14365 30035 14399
rect 3985 14297 4019 14331
rect 6469 14297 6503 14331
rect 11630 14297 11664 14331
rect 12725 14297 12759 14331
rect 25973 14297 26007 14331
rect 28825 14297 28859 14331
rect 2973 14229 3007 14263
rect 4185 14229 4219 14263
rect 4353 14229 4387 14263
rect 7389 14229 7423 14263
rect 9597 14229 9631 14263
rect 12541 14229 12575 14263
rect 15669 14229 15703 14263
rect 16313 14229 16347 14263
rect 18245 14229 18279 14263
rect 26249 14229 26283 14263
rect 28089 14229 28123 14263
rect 31125 14229 31159 14263
rect 10609 14025 10643 14059
rect 11713 14025 11747 14059
rect 13277 14025 13311 14059
rect 14105 14025 14139 14059
rect 16221 14025 16255 14059
rect 18429 14025 18463 14059
rect 5641 13957 5675 13991
rect 5857 13957 5891 13991
rect 8217 13957 8251 13991
rect 15301 13957 15335 13991
rect 15853 13957 15887 13991
rect 19717 13957 19751 13991
rect 30297 13957 30331 13991
rect 30497 13957 30531 13991
rect 1777 13889 1811 13923
rect 1961 13889 1995 13923
rect 2605 13889 2639 13923
rect 3249 13889 3283 13923
rect 3433 13889 3467 13923
rect 3525 13889 3559 13923
rect 3617 13889 3651 13923
rect 4537 13889 4571 13923
rect 7021 13889 7055 13923
rect 9229 13889 9263 13923
rect 9485 13889 9519 13923
rect 11897 13889 11931 13923
rect 13553 13889 13587 13923
rect 14289 13889 14323 13923
rect 15025 13889 15059 13923
rect 15761 13889 15795 13923
rect 16037 13889 16071 13923
rect 17325 13889 17359 13923
rect 22017 13889 22051 13923
rect 22477 13889 22511 13923
rect 23213 13889 23247 13923
rect 23305 13889 23339 13923
rect 24225 13889 24259 13923
rect 24501 13889 24535 13923
rect 25237 13889 25271 13923
rect 25697 13889 25731 13923
rect 26433 13889 26467 13923
rect 26525 13889 26559 13923
rect 27721 13889 27755 13923
rect 27977 13889 28011 13923
rect 29561 13889 29595 13923
rect 29745 13889 29779 13923
rect 29837 13889 29871 13923
rect 31125 13889 31159 13923
rect 2789 13821 2823 13855
rect 3893 13821 3927 13855
rect 4445 13821 4479 13855
rect 13277 13821 13311 13855
rect 13461 13821 13495 13855
rect 15117 13821 15151 13855
rect 22293 13821 22327 13855
rect 25513 13821 25547 13855
rect 6745 13753 6779 13787
rect 24409 13753 24443 13787
rect 29561 13753 29595 13787
rect 30665 13753 30699 13787
rect 31309 13753 31343 13787
rect 1961 13685 1995 13719
rect 2421 13685 2455 13719
rect 4813 13685 4847 13719
rect 5825 13685 5859 13719
rect 6009 13685 6043 13719
rect 6561 13685 6595 13719
rect 8125 13685 8159 13719
rect 14841 13685 14875 13719
rect 15301 13685 15335 13719
rect 17509 13685 17543 13719
rect 22477 13685 22511 13719
rect 22661 13685 22695 13719
rect 24317 13685 24351 13719
rect 25329 13685 25363 13719
rect 25881 13685 25915 13719
rect 29101 13685 29135 13719
rect 30481 13685 30515 13719
rect 4169 13481 4203 13515
rect 5365 13481 5399 13515
rect 7113 13481 7147 13515
rect 10425 13481 10459 13515
rect 10609 13481 10643 13515
rect 18797 13481 18831 13515
rect 22109 13481 22143 13515
rect 25973 13481 26007 13515
rect 27813 13481 27847 13515
rect 28365 13481 28399 13515
rect 3433 13413 3467 13447
rect 4353 13413 4387 13447
rect 9505 13413 9539 13447
rect 12909 13413 12943 13447
rect 19441 13413 19475 13447
rect 21925 13413 21959 13447
rect 25605 13413 25639 13447
rect 26801 13413 26835 13447
rect 29193 13413 29227 13447
rect 5181 13345 5215 13379
rect 6009 13345 6043 13379
rect 6101 13345 6135 13379
rect 14565 13345 14599 13379
rect 14657 13345 14691 13379
rect 20177 13345 20211 13379
rect 22293 13345 22327 13379
rect 23489 13345 23523 13379
rect 25973 13345 26007 13379
rect 27721 13345 27755 13379
rect 30205 13345 30239 13379
rect 2237 13277 2271 13311
rect 2697 13277 2731 13311
rect 2881 13277 2915 13311
rect 2973 13277 3007 13311
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 4905 13277 4939 13311
rect 5365 13277 5399 13311
rect 6377 13277 6411 13311
rect 6469 13277 6503 13311
rect 7297 13277 7331 13311
rect 7389 13277 7423 13311
rect 7573 13277 7607 13311
rect 7665 13277 7699 13311
rect 9505 13277 9539 13311
rect 9781 13277 9815 13311
rect 11253 13277 11287 13311
rect 11989 13277 12023 13311
rect 12173 13277 12207 13311
rect 12909 13277 12943 13311
rect 13093 13277 13127 13311
rect 13737 13277 13771 13311
rect 14473 13277 14507 13311
rect 14749 13277 14783 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 17417 13277 17451 13311
rect 17673 13277 17707 13311
rect 19717 13277 19751 13311
rect 20361 13277 20395 13311
rect 20453 13277 20487 13311
rect 21465 13277 21499 13311
rect 22109 13277 22143 13311
rect 23397 13277 23431 13311
rect 24593 13277 24627 13311
rect 24777 13277 24811 13311
rect 25789 13277 25823 13311
rect 26709 13277 26743 13311
rect 27629 13277 27663 13311
rect 28273 13277 28307 13311
rect 28457 13277 28491 13311
rect 28917 13277 28951 13311
rect 29193 13277 29227 13311
rect 30021 13277 30055 13311
rect 3985 13209 4019 13243
rect 4185 13209 4219 13243
rect 10577 13209 10611 13243
rect 10793 13209 10827 13243
rect 19441 13209 19475 13243
rect 20177 13209 20211 13243
rect 22569 13209 22603 13243
rect 24685 13209 24719 13243
rect 26249 13209 26283 13243
rect 27353 13209 27387 13243
rect 29745 13209 29779 13243
rect 2145 13141 2179 13175
rect 5549 13141 5583 13175
rect 6285 13141 6319 13175
rect 6653 13141 6687 13175
rect 9689 13141 9723 13175
rect 11437 13141 11471 13175
rect 12081 13141 12115 13175
rect 13553 13141 13587 13175
rect 14289 13141 14323 13175
rect 15393 13141 15427 13175
rect 19625 13141 19659 13175
rect 21373 13141 21407 13175
rect 23029 13141 23063 13175
rect 27445 13141 27479 13175
rect 29009 13141 29043 13175
rect 29837 13141 29871 13175
rect 2881 12937 2915 12971
rect 4905 12937 4939 12971
rect 5825 12937 5859 12971
rect 5917 12937 5951 12971
rect 8125 12937 8159 12971
rect 9321 12937 9355 12971
rect 18337 12937 18371 12971
rect 22017 12937 22051 12971
rect 22661 12937 22695 12971
rect 23673 12937 23707 12971
rect 24685 12937 24719 12971
rect 26341 12937 26375 12971
rect 27445 12937 27479 12971
rect 2329 12869 2363 12903
rect 4137 12869 4171 12903
rect 4353 12869 4387 12903
rect 5733 12869 5767 12903
rect 15393 12869 15427 12903
rect 19450 12869 19484 12903
rect 25973 12869 26007 12903
rect 28273 12869 28307 12903
rect 28457 12869 28491 12903
rect 2237 12801 2271 12835
rect 2421 12801 2455 12835
rect 3065 12801 3099 12835
rect 3157 12801 3191 12835
rect 3249 12801 3283 12835
rect 3341 12801 3375 12835
rect 3525 12801 3559 12835
rect 4813 12801 4847 12835
rect 4997 12801 5031 12835
rect 5641 12801 5675 12835
rect 6009 12801 6043 12835
rect 7012 12801 7046 12835
rect 9505 12801 9539 12835
rect 9689 12801 9723 12835
rect 10517 12801 10551 12835
rect 13185 12801 13219 12835
rect 13452 12801 13486 12835
rect 15025 12801 15059 12835
rect 15209 12801 15243 12835
rect 15301 12801 15335 12835
rect 15531 12801 15565 12835
rect 21189 12801 21223 12835
rect 22293 12801 22327 12835
rect 22753 12801 22787 12835
rect 23305 12801 23339 12835
rect 23732 12801 23766 12835
rect 24317 12801 24351 12835
rect 24501 12801 24535 12835
rect 25697 12801 25731 12835
rect 25790 12801 25824 12835
rect 26065 12801 26099 12835
rect 26162 12801 26196 12835
rect 27353 12801 27387 12835
rect 27629 12801 27663 12835
rect 28641 12801 28675 12835
rect 29101 12801 29135 12835
rect 29377 12801 29411 12835
rect 29653 12801 29687 12835
rect 29837 12801 29871 12835
rect 30564 12801 30598 12835
rect 6745 12733 6779 12767
rect 10609 12733 10643 12767
rect 15669 12733 15703 12767
rect 19717 12733 19751 12767
rect 21465 12733 21499 12767
rect 23213 12733 23247 12767
rect 29469 12733 29503 12767
rect 30297 12733 30331 12767
rect 14565 12665 14599 12699
rect 21281 12665 21315 12699
rect 21373 12665 21407 12699
rect 22477 12665 22511 12699
rect 23857 12665 23891 12699
rect 27629 12665 27663 12699
rect 29561 12665 29595 12699
rect 3985 12597 4019 12631
rect 4169 12597 4203 12631
rect 10241 12597 10275 12631
rect 22385 12597 22419 12631
rect 31677 12597 31711 12631
rect 4169 12393 4203 12427
rect 6377 12393 6411 12427
rect 7021 12393 7055 12427
rect 9689 12393 9723 12427
rect 11529 12393 11563 12427
rect 13553 12393 13587 12427
rect 13737 12393 13771 12427
rect 15485 12393 15519 12427
rect 15669 12393 15703 12427
rect 21557 12393 21591 12427
rect 22017 12393 22051 12427
rect 23213 12393 23247 12427
rect 26341 12393 26375 12427
rect 27721 12393 27755 12427
rect 30757 12393 30791 12427
rect 2973 12325 3007 12359
rect 14289 12325 14323 12359
rect 28365 12325 28399 12359
rect 2513 12257 2547 12291
rect 4261 12257 4295 12291
rect 9413 12257 9447 12291
rect 17141 12257 17175 12291
rect 21281 12257 21315 12291
rect 22477 12257 22511 12291
rect 22569 12257 22603 12291
rect 25973 12257 26007 12291
rect 30021 12257 30055 12291
rect 30113 12257 30147 12291
rect 2605 12189 2639 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 7205 12189 7239 12223
rect 9321 12189 9355 12223
rect 10149 12189 10183 12223
rect 12081 12189 12115 12223
rect 12357 12189 12391 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 14841 12189 14875 12223
rect 17233 12189 17267 12223
rect 18245 12189 18279 12223
rect 18521 12189 18555 12223
rect 21189 12189 21223 12223
rect 23213 12189 23247 12223
rect 23397 12189 23431 12223
rect 24777 12189 24811 12223
rect 24961 12189 24995 12223
rect 25605 12189 25639 12223
rect 25789 12189 25823 12223
rect 25881 12189 25915 12223
rect 26157 12189 26191 12223
rect 27997 12189 28031 12223
rect 28457 12189 28491 12223
rect 29101 12189 29135 12223
rect 29193 12189 29227 12223
rect 29929 12189 29963 12223
rect 30205 12189 30239 12223
rect 30941 12189 30975 12223
rect 6361 12121 6395 12155
rect 6561 12121 6595 12155
rect 10416 12121 10450 12155
rect 13369 12121 13403 12155
rect 14657 12121 14691 12155
rect 15301 12121 15335 12155
rect 18061 12121 18095 12155
rect 18429 12121 18463 12155
rect 22385 12121 22419 12155
rect 28917 12121 28951 12155
rect 6193 12053 6227 12087
rect 12173 12053 12207 12087
rect 12541 12053 12575 12087
rect 13579 12053 13613 12087
rect 15511 12053 15545 12087
rect 17601 12053 17635 12087
rect 25145 12053 25179 12087
rect 28089 12053 28123 12087
rect 28181 12053 28215 12087
rect 29015 12053 29049 12087
rect 29745 12053 29779 12087
rect 3065 11849 3099 11883
rect 18613 11849 18647 11883
rect 26433 11849 26467 11883
rect 28181 11849 28215 11883
rect 29377 11849 29411 11883
rect 29929 11849 29963 11883
rect 10916 11781 10950 11815
rect 14657 11781 14691 11815
rect 16957 11781 16991 11815
rect 18153 11781 18187 11815
rect 3249 11713 3283 11747
rect 4885 11713 4919 11747
rect 6745 11713 6779 11747
rect 6929 11713 6963 11747
rect 11161 11713 11195 11747
rect 13645 11713 13679 11747
rect 14473 11713 14507 11747
rect 15393 11713 15427 11747
rect 16313 11713 16347 11747
rect 16865 11713 16899 11747
rect 17049 11713 17083 11747
rect 17785 11713 17819 11747
rect 18797 11713 18831 11747
rect 19073 11713 19107 11747
rect 22385 11713 22419 11747
rect 23581 11713 23615 11747
rect 23765 11713 23799 11747
rect 26525 11713 26559 11747
rect 27169 11713 27203 11747
rect 27905 11713 27939 11747
rect 27997 11713 28031 11747
rect 28733 11713 28767 11747
rect 28917 11713 28951 11747
rect 29009 11713 29043 11747
rect 29101 11713 29135 11747
rect 29837 11713 29871 11747
rect 30021 11713 30055 11747
rect 30665 11713 30699 11747
rect 3433 11645 3467 11679
rect 4629 11645 4663 11679
rect 7021 11645 7055 11679
rect 15121 11645 15155 11679
rect 15301 11645 15335 11679
rect 16221 11645 16255 11679
rect 17693 11645 17727 11679
rect 18061 11645 18095 11679
rect 18889 11645 18923 11679
rect 22477 11645 22511 11679
rect 27445 11645 27479 11679
rect 28181 11645 28215 11679
rect 30573 11645 30607 11679
rect 17509 11577 17543 11611
rect 22017 11577 22051 11611
rect 27261 11577 27295 11611
rect 6009 11509 6043 11543
rect 6561 11509 6595 11543
rect 9781 11509 9815 11543
rect 13461 11509 13495 11543
rect 14381 11509 14415 11543
rect 15209 11509 15243 11543
rect 15945 11509 15979 11543
rect 16313 11509 16347 11543
rect 19073 11509 19107 11543
rect 23673 11509 23707 11543
rect 27353 11509 27387 11543
rect 30941 11509 30975 11543
rect 4905 11305 4939 11339
rect 5733 11305 5767 11339
rect 9781 11305 9815 11339
rect 10425 11305 10459 11339
rect 16865 11305 16899 11339
rect 17509 11305 17543 11339
rect 19441 11305 19475 11339
rect 25145 11305 25179 11339
rect 29837 11305 29871 11339
rect 30205 11305 30239 11339
rect 30757 11305 30791 11339
rect 30941 11305 30975 11339
rect 4261 11237 4295 11271
rect 6561 11237 6595 11271
rect 6929 11237 6963 11271
rect 16681 11237 16715 11271
rect 20177 11237 20211 11271
rect 22569 11237 22603 11271
rect 26801 11237 26835 11271
rect 28181 11237 28215 11271
rect 29101 11237 29135 11271
rect 2973 11169 3007 11203
rect 15485 11169 15519 11203
rect 18153 11169 18187 11203
rect 19717 11169 19751 11203
rect 20729 11169 20763 11203
rect 21005 11169 21039 11203
rect 23581 11169 23615 11203
rect 24685 11169 24719 11203
rect 27629 11169 27663 11203
rect 31033 11169 31067 11203
rect 2881 11101 2915 11135
rect 3985 11101 4019 11135
rect 4905 11101 4939 11135
rect 5089 11101 5123 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 6745 11101 6779 11135
rect 7757 11101 7791 11135
rect 8401 11101 8435 11135
rect 9689 11101 9723 11135
rect 9873 11101 9907 11135
rect 10425 11101 10459 11135
rect 10609 11101 10643 11135
rect 14289 11101 14323 11135
rect 14565 11101 14599 11135
rect 15393 11101 15427 11135
rect 17693 11101 17727 11135
rect 17785 11101 17819 11135
rect 21097 11101 21131 11135
rect 22753 11101 22787 11135
rect 22845 11101 22879 11135
rect 23121 11101 23155 11135
rect 23765 11101 23799 11135
rect 23949 11101 23983 11135
rect 24777 11101 24811 11135
rect 25789 11101 25823 11135
rect 25881 11101 25915 11135
rect 26525 11101 26559 11135
rect 27997 11101 28031 11135
rect 28917 11101 28951 11135
rect 29193 11101 29227 11135
rect 29745 11101 29779 11135
rect 31309 11101 31343 11135
rect 4261 11033 4295 11067
rect 5717 11033 5751 11067
rect 5917 11033 5951 11067
rect 7389 11033 7423 11067
rect 14749 11033 14783 11067
rect 16833 11033 16867 11067
rect 17049 11033 17083 11067
rect 18061 11033 18095 11067
rect 20177 11033 20211 11067
rect 22937 11033 22971 11067
rect 26801 11033 26835 11067
rect 27905 11033 27939 11067
rect 2513 10965 2547 10999
rect 4077 10965 4111 10999
rect 5549 10965 5583 10999
rect 8585 10965 8619 10999
rect 14381 10965 14415 10999
rect 15761 10965 15795 10999
rect 19625 10965 19659 10999
rect 26065 10965 26099 10999
rect 26617 10965 26651 10999
rect 27813 10965 27847 10999
rect 28733 10965 28767 10999
rect 2605 10761 2639 10795
rect 3617 10761 3651 10795
rect 10057 10761 10091 10795
rect 15853 10761 15887 10795
rect 17417 10761 17451 10795
rect 18153 10761 18187 10795
rect 19809 10761 19843 10795
rect 25605 10761 25639 10795
rect 31309 10761 31343 10795
rect 9597 10693 9631 10727
rect 13001 10693 13035 10727
rect 14749 10693 14783 10727
rect 19165 10693 19199 10727
rect 23397 10693 23431 10727
rect 30481 10693 30515 10727
rect 2329 10625 2363 10659
rect 3157 10625 3191 10659
rect 3433 10625 3467 10659
rect 5365 10625 5399 10659
rect 5825 10625 5859 10659
rect 10241 10625 10275 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 15209 10625 15243 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 15577 10625 15611 10659
rect 15669 10625 15703 10659
rect 17049 10625 17083 10659
rect 18337 10625 18371 10659
rect 18429 10625 18463 10659
rect 18613 10625 18647 10659
rect 18705 10625 18739 10659
rect 19625 10625 19659 10659
rect 20637 10625 20671 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 22293 10625 22327 10659
rect 22385 10625 22419 10659
rect 25973 10625 26007 10659
rect 27537 10625 27571 10659
rect 27721 10625 27755 10659
rect 28733 10625 28767 10659
rect 28917 10625 28951 10659
rect 29837 10625 29871 10659
rect 30021 10625 30055 10659
rect 30665 10625 30699 10659
rect 30757 10625 30791 10659
rect 31217 10625 31251 10659
rect 31493 10625 31527 10659
rect 2605 10557 2639 10591
rect 3341 10557 3375 10591
rect 10425 10557 10459 10591
rect 17141 10557 17175 10591
rect 19441 10557 19475 10591
rect 20545 10557 20579 10591
rect 26065 10557 26099 10591
rect 28825 10557 28859 10591
rect 29009 10557 29043 10591
rect 2421 10489 2455 10523
rect 3249 10489 3283 10523
rect 29193 10489 29227 10523
rect 30481 10489 30515 10523
rect 5181 10421 5215 10455
rect 6009 10421 6043 10455
rect 8309 10421 8343 10455
rect 11713 10421 11747 10455
rect 19625 10421 19659 10455
rect 20361 10421 20395 10455
rect 22661 10421 22695 10455
rect 24685 10421 24719 10455
rect 27905 10421 27939 10455
rect 29653 10421 29687 10455
rect 29837 10421 29871 10455
rect 31493 10421 31527 10455
rect 2697 10217 2731 10251
rect 3065 10217 3099 10251
rect 3157 10217 3191 10251
rect 7941 10217 7975 10251
rect 10517 10217 10551 10251
rect 14289 10217 14323 10251
rect 17509 10217 17543 10251
rect 18705 10217 18739 10251
rect 19993 10217 20027 10251
rect 23029 10217 23063 10251
rect 23949 10217 23983 10251
rect 27629 10217 27663 10251
rect 31033 10217 31067 10251
rect 31769 10217 31803 10251
rect 3249 10149 3283 10183
rect 15117 10149 15151 10183
rect 18521 10149 18555 10183
rect 19441 10149 19475 10183
rect 14473 10081 14507 10115
rect 14657 10081 14691 10115
rect 16589 10081 16623 10115
rect 20913 10081 20947 10115
rect 25513 10081 25547 10115
rect 27169 10081 27203 10115
rect 28457 10081 28491 10115
rect 28549 10081 28583 10115
rect 30205 10081 30239 10115
rect 30941 10081 30975 10115
rect 2053 10013 2087 10047
rect 2237 10013 2271 10047
rect 2973 10013 3007 10047
rect 3433 10013 3467 10047
rect 4629 10013 4663 10047
rect 6561 10013 6595 10047
rect 9137 10013 9171 10047
rect 11069 10013 11103 10047
rect 12909 10013 12943 10047
rect 14565 10013 14599 10047
rect 15301 10013 15335 10047
rect 15577 10013 15611 10047
rect 16497 10013 16531 10047
rect 19625 10013 19659 10047
rect 22569 10013 22603 10047
rect 23857 10013 23891 10047
rect 24041 10013 24075 10047
rect 24994 10013 25028 10047
rect 25421 10013 25455 10047
rect 26157 10013 26191 10047
rect 26341 10013 26375 10047
rect 26525 10013 26559 10047
rect 27353 10013 27387 10047
rect 27445 10013 27479 10047
rect 27721 10013 27755 10047
rect 28365 10013 28399 10047
rect 28641 10013 28675 10047
rect 30113 10013 30147 10047
rect 31125 10013 31159 10047
rect 31309 10013 31343 10047
rect 31769 10013 31803 10047
rect 31953 10013 31987 10047
rect 2145 9945 2179 9979
rect 4896 9945 4930 9979
rect 6828 9945 6862 9979
rect 9382 9945 9416 9979
rect 11336 9945 11370 9979
rect 13001 9945 13035 9979
rect 13185 9945 13219 9979
rect 14289 9945 14323 9979
rect 17693 9945 17727 9979
rect 18889 9945 18923 9979
rect 19717 9945 19751 9979
rect 23213 9945 23247 9979
rect 23397 9945 23431 9979
rect 26249 9945 26283 9979
rect 30849 9945 30883 9979
rect 6009 9877 6043 9911
rect 12449 9877 12483 9911
rect 12909 9877 12943 9911
rect 15485 9877 15519 9911
rect 16865 9877 16899 9911
rect 17325 9877 17359 9911
rect 17493 9877 17527 9911
rect 18679 9877 18713 9911
rect 19809 9877 19843 9911
rect 24869 9877 24903 9911
rect 25053 9877 25087 9911
rect 25973 9877 26007 9911
rect 28181 9877 28215 9911
rect 29745 9877 29779 9911
rect 30389 9877 30423 9911
rect 1961 9673 1995 9707
rect 2421 9673 2455 9707
rect 14381 9673 14415 9707
rect 20453 9673 20487 9707
rect 22201 9673 22235 9707
rect 25421 9673 25455 9707
rect 27905 9673 27939 9707
rect 31677 9673 31711 9707
rect 1593 9605 1627 9639
rect 1809 9605 1843 9639
rect 3433 9605 3467 9639
rect 4353 9605 4387 9639
rect 6009 9605 6043 9639
rect 9321 9605 9355 9639
rect 9537 9605 9571 9639
rect 15209 9605 15243 9639
rect 16313 9605 16347 9639
rect 18613 9605 18647 9639
rect 25329 9605 25363 9639
rect 26249 9605 26283 9639
rect 26465 9605 26499 9639
rect 28917 9605 28951 9639
rect 30564 9605 30598 9639
rect 2789 9537 2823 9571
rect 3709 9537 3743 9571
rect 4169 9537 4203 9571
rect 4445 9537 4479 9571
rect 4537 9537 4571 9571
rect 5825 9537 5859 9571
rect 6929 9537 6963 9571
rect 7185 9537 7219 9571
rect 10149 9537 10183 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 10517 9537 10551 9571
rect 11897 9537 11931 9571
rect 12081 9537 12115 9571
rect 12173 9537 12207 9571
rect 13001 9537 13035 9571
rect 13268 9537 13302 9571
rect 15025 9537 15059 9571
rect 15301 9537 15335 9571
rect 16129 9537 16163 9571
rect 18337 9537 18371 9571
rect 19257 9537 19291 9571
rect 19441 9537 19475 9571
rect 19533 9537 19567 9571
rect 20821 9537 20855 9571
rect 22017 9537 22051 9571
rect 22201 9537 22235 9571
rect 22928 9537 22962 9571
rect 27537 9537 27571 9571
rect 27629 9537 27663 9571
rect 28549 9537 28583 9571
rect 28733 9537 28767 9571
rect 29377 9537 29411 9571
rect 29469 9537 29503 9571
rect 30297 9537 30331 9571
rect 2697 9469 2731 9503
rect 3433 9469 3467 9503
rect 5641 9469 5675 9503
rect 10793 9469 10827 9503
rect 15945 9469 15979 9503
rect 18613 9469 18647 9503
rect 19073 9469 19107 9503
rect 20729 9469 20763 9503
rect 22661 9469 22695 9503
rect 25605 9469 25639 9503
rect 29653 9469 29687 9503
rect 11713 9401 11747 9435
rect 18429 9401 18463 9435
rect 24041 9401 24075 9435
rect 1777 9333 1811 9367
rect 3617 9333 3651 9367
rect 4721 9333 4755 9367
rect 8309 9333 8343 9367
rect 9505 9333 9539 9367
rect 9689 9333 9723 9367
rect 14841 9333 14875 9367
rect 24961 9333 24995 9367
rect 26433 9333 26467 9367
rect 26617 9333 26651 9367
rect 27721 9333 27755 9367
rect 29561 9333 29595 9367
rect 3433 9129 3467 9163
rect 5825 9129 5859 9163
rect 6561 9129 6595 9163
rect 10057 9129 10091 9163
rect 13001 9129 13035 9163
rect 18705 9129 18739 9163
rect 20821 9129 20855 9163
rect 26617 9129 26651 9163
rect 27077 9129 27111 9163
rect 29837 9129 29871 9163
rect 2421 9061 2455 9095
rect 3157 9061 3191 9095
rect 8493 9061 8527 9095
rect 10701 9061 10735 9095
rect 15853 9061 15887 9095
rect 27629 9061 27663 9095
rect 28917 9061 28951 9095
rect 1961 8993 1995 9027
rect 3065 8993 3099 9027
rect 6929 8993 6963 9027
rect 14473 8993 14507 9027
rect 24593 8993 24627 9027
rect 28089 8993 28123 9027
rect 28181 8993 28215 9027
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 6745 8925 6779 8959
rect 7389 8925 7423 8959
rect 7757 8925 7791 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 9505 8925 9539 8959
rect 9873 8925 9907 8959
rect 11814 8925 11848 8959
rect 12081 8925 12115 8959
rect 12817 8925 12851 8959
rect 13553 8925 13587 8959
rect 13737 8925 13771 8959
rect 14740 8925 14774 8959
rect 16313 8925 16347 8959
rect 16497 8925 16531 8959
rect 19441 8925 19475 8959
rect 21281 8925 21315 8959
rect 21465 8925 21499 8959
rect 22201 8925 22235 8959
rect 22468 8925 22502 8959
rect 24777 8925 24811 8959
rect 25881 8925 25915 8959
rect 25973 8925 26007 8959
rect 26801 8925 26835 8959
rect 26893 8925 26927 8959
rect 27169 8925 27203 8959
rect 27997 8925 28031 8959
rect 28825 8925 28859 8959
rect 29009 8925 29043 8959
rect 29745 8925 29779 8959
rect 29929 8925 29963 8959
rect 30573 8925 30607 8959
rect 5457 8857 5491 8891
rect 5641 8857 5675 8891
rect 7573 8857 7607 8891
rect 7665 8857 7699 8891
rect 9689 8857 9723 8891
rect 9781 8857 9815 8891
rect 12633 8857 12667 8891
rect 13645 8857 13679 8891
rect 18521 8857 18555 8891
rect 19708 8857 19742 8891
rect 26157 8857 26191 8891
rect 7941 8789 7975 8823
rect 16313 8789 16347 8823
rect 18721 8789 18755 8823
rect 18889 8789 18923 8823
rect 23581 8789 23615 8823
rect 24961 8789 24995 8823
rect 30389 8789 30423 8823
rect 2973 8585 3007 8619
rect 5457 8585 5491 8619
rect 7757 8585 7791 8619
rect 9873 8585 9907 8619
rect 10977 8585 11011 8619
rect 12633 8585 12667 8619
rect 14933 8585 14967 8619
rect 18613 8585 18647 8619
rect 19901 8585 19935 8619
rect 22385 8585 22419 8619
rect 24317 8585 24351 8619
rect 26525 8585 26559 8619
rect 30941 8585 30975 8619
rect 3433 8517 3467 8551
rect 11713 8517 11747 8551
rect 1777 8449 1811 8483
rect 1961 8449 1995 8483
rect 2605 8449 2639 8483
rect 3617 8449 3651 8483
rect 5641 8449 5675 8483
rect 5733 8449 5767 8483
rect 6009 8449 6043 8483
rect 6561 8449 6595 8483
rect 7849 8449 7883 8483
rect 8585 8449 8619 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 10517 8449 10551 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 12541 8449 12575 8483
rect 12725 8449 12759 8483
rect 13277 8449 13311 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 14197 8449 14231 8483
rect 16057 8449 16091 8483
rect 16313 8449 16347 8483
rect 17233 8449 17267 8483
rect 17500 8449 17534 8483
rect 21025 8449 21059 8483
rect 21281 8449 21315 8483
rect 23498 8449 23532 8483
rect 23765 8449 23799 8483
rect 24225 8449 24259 8483
rect 24409 8449 24443 8483
rect 25145 8449 25179 8483
rect 25412 8449 25446 8483
rect 27169 8449 27203 8483
rect 27425 8449 27459 8483
rect 29561 8449 29595 8483
rect 29828 8449 29862 8483
rect 1869 8381 1903 8415
rect 2513 8381 2547 8415
rect 3893 8381 3927 8415
rect 5917 8381 5951 8415
rect 8769 8381 8803 8415
rect 10609 8381 10643 8415
rect 3801 8313 3835 8347
rect 8401 8313 8435 8347
rect 11713 8313 11747 8347
rect 13461 8313 13495 8347
rect 6745 8245 6779 8279
rect 10333 8245 10367 8279
rect 28549 8245 28583 8279
rect 2789 8041 2823 8075
rect 6745 8041 6779 8075
rect 8585 8041 8619 8075
rect 9321 8041 9355 8075
rect 16957 8041 16991 8075
rect 17601 8041 17635 8075
rect 19901 8041 19935 8075
rect 21189 8041 21223 8075
rect 23673 8041 23707 8075
rect 25421 8041 25455 8075
rect 26985 8041 27019 8075
rect 27997 8041 28031 8075
rect 10241 7973 10275 8007
rect 20729 7973 20763 8007
rect 23029 7973 23063 8007
rect 24593 7973 24627 8007
rect 5917 7905 5951 7939
rect 7205 7905 7239 7939
rect 14473 7905 14507 7939
rect 16773 7905 16807 7939
rect 19441 7905 19475 7939
rect 27721 7905 27755 7939
rect 2789 7837 2823 7871
rect 2973 7837 3007 7871
rect 6561 7837 6595 7871
rect 9965 7837 9999 7871
rect 11161 7837 11195 7871
rect 11345 7837 11379 7871
rect 11805 7837 11839 7871
rect 14729 7837 14763 7871
rect 16681 7837 16715 7871
rect 17417 7837 17451 7871
rect 17601 7837 17635 7871
rect 19533 7837 19567 7871
rect 19717 7837 19751 7871
rect 20453 7837 20487 7871
rect 21189 7837 21223 7871
rect 21373 7837 21407 7871
rect 22753 7837 22787 7871
rect 22845 7837 22879 7871
rect 24593 7837 24627 7871
rect 24777 7837 24811 7871
rect 25237 7837 25271 7871
rect 26801 7837 26835 7871
rect 27629 7837 27663 7871
rect 5672 7769 5706 7803
rect 7450 7769 7484 7803
rect 9305 7769 9339 7803
rect 9505 7769 9539 7803
rect 10241 7769 10275 7803
rect 11253 7769 11287 7803
rect 12050 7769 12084 7803
rect 16313 7769 16347 7803
rect 16405 7769 16439 7803
rect 20729 7769 20763 7803
rect 23029 7769 23063 7803
rect 23857 7769 23891 7803
rect 4537 7701 4571 7735
rect 9137 7701 9171 7735
rect 10057 7701 10091 7735
rect 13185 7701 13219 7735
rect 15853 7701 15887 7735
rect 20545 7701 20579 7735
rect 23489 7701 23523 7735
rect 23657 7701 23691 7735
rect 2881 7497 2915 7531
rect 3065 7497 3099 7531
rect 4445 7497 4479 7531
rect 5825 7497 5859 7531
rect 6837 7497 6871 7531
rect 9137 7497 9171 7531
rect 9505 7497 9539 7531
rect 12173 7497 12207 7531
rect 12357 7497 12391 7531
rect 14105 7497 14139 7531
rect 15393 7497 15427 7531
rect 16313 7497 16347 7531
rect 17693 7497 17727 7531
rect 17877 7497 17911 7531
rect 19993 7497 20027 7531
rect 20161 7497 20195 7531
rect 22753 7497 22787 7531
rect 23857 7497 23891 7531
rect 24317 7497 24351 7531
rect 25237 7497 25271 7531
rect 7665 7429 7699 7463
rect 9965 7429 9999 7463
rect 10165 7429 10199 7463
rect 11069 7429 11103 7463
rect 20361 7429 20395 7463
rect 24685 7429 24719 7463
rect 25329 7429 25363 7463
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 4077 7361 4111 7395
rect 5457 7361 5491 7395
rect 5828 7361 5862 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 7389 7361 7423 7395
rect 7481 7361 7515 7395
rect 8125 7361 8159 7395
rect 8401 7361 8435 7395
rect 9045 7361 9079 7395
rect 9321 7361 9355 7395
rect 10793 7361 10827 7395
rect 10885 7361 10919 7395
rect 12298 7361 12332 7395
rect 13553 7361 13587 7395
rect 13737 7361 13771 7395
rect 13829 7361 13863 7395
rect 13921 7361 13955 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 16129 7361 16163 7395
rect 17752 7361 17786 7395
rect 22569 7361 22603 7395
rect 22753 7361 22787 7395
rect 23397 7361 23431 7395
rect 24501 7361 24535 7395
rect 24777 7361 24811 7395
rect 25237 7361 25271 7395
rect 25513 7361 25547 7395
rect 4169 7293 4203 7327
rect 5365 7293 5399 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 15853 7293 15887 7327
rect 17233 7293 17267 7327
rect 17325 7293 17359 7327
rect 20821 7293 20855 7327
rect 23489 7293 23523 7327
rect 3433 7225 3467 7259
rect 7665 7225 7699 7259
rect 8217 7225 8251 7259
rect 10793 7225 10827 7259
rect 21097 7225 21131 7259
rect 23213 7225 23247 7259
rect 2329 7157 2363 7191
rect 3065 7157 3099 7191
rect 6009 7157 6043 7191
rect 8585 7157 8619 7191
rect 10149 7157 10183 7191
rect 10333 7157 10367 7191
rect 15945 7157 15979 7191
rect 20177 7157 20211 7191
rect 21281 7157 21315 7191
rect 4169 6953 4203 6987
rect 5273 6953 5307 6987
rect 5917 6953 5951 6987
rect 6561 6953 6595 6987
rect 13093 6953 13127 6987
rect 16037 6953 16071 6987
rect 17417 6953 17451 6987
rect 17969 6953 18003 6987
rect 20453 6953 20487 6987
rect 22569 6953 22603 6987
rect 23857 6953 23891 6987
rect 3065 6885 3099 6919
rect 12541 6885 12575 6919
rect 14381 6885 14415 6919
rect 22385 6885 22419 6919
rect 2605 6817 2639 6851
rect 4997 6817 5031 6851
rect 7665 6817 7699 6851
rect 9321 6817 9355 6851
rect 9413 6817 9447 6851
rect 10333 6817 10367 6851
rect 12265 6817 12299 6851
rect 13277 6817 13311 6851
rect 14749 6817 14783 6851
rect 17141 6817 17175 6851
rect 21925 6817 21959 6851
rect 2743 6749 2777 6783
rect 4077 6749 4111 6783
rect 4261 6749 4295 6783
rect 4905 6749 4939 6783
rect 5733 6749 5767 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 7573 6749 7607 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 9781 6749 9815 6783
rect 10241 6749 10275 6783
rect 10425 6749 10459 6783
rect 11253 6749 11287 6783
rect 11529 6749 11563 6783
rect 12173 6749 12207 6783
rect 13369 6749 13403 6783
rect 15945 6749 15979 6783
rect 17049 6749 17083 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 19441 6749 19475 6783
rect 20637 6749 20671 6783
rect 20729 6749 20763 6783
rect 20913 6749 20947 6783
rect 21005 6749 21039 6783
rect 21465 6749 21499 6783
rect 21557 6749 21591 6783
rect 21741 6749 21775 6783
rect 23673 6749 23707 6783
rect 8585 6681 8619 6715
rect 11069 6681 11103 6715
rect 22537 6681 22571 6715
rect 22753 6681 22787 6715
rect 23489 6681 23523 6715
rect 9137 6613 9171 6647
rect 9597 6613 9631 6647
rect 9689 6613 9723 6647
rect 11437 6613 11471 6647
rect 14289 6613 14323 6647
rect 16405 6613 16439 6647
rect 19625 6613 19659 6647
rect 4261 6409 4295 6443
rect 9505 6409 9539 6443
rect 13461 6409 13495 6443
rect 16865 6409 16899 6443
rect 20085 6409 20119 6443
rect 22017 6409 22051 6443
rect 4353 6341 4387 6375
rect 4905 6341 4939 6375
rect 5089 6341 5123 6375
rect 5273 6341 5307 6375
rect 7941 6341 7975 6375
rect 19625 6341 19659 6375
rect 3985 6273 4019 6307
rect 4445 6273 4479 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 8493 6273 8527 6307
rect 8677 6273 8711 6307
rect 9321 6273 9355 6307
rect 9505 6273 9539 6307
rect 11989 6273 12023 6307
rect 13093 6273 13127 6307
rect 14749 6273 14783 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 16129 6273 16163 6307
rect 17049 6273 17083 6307
rect 18429 6273 18463 6307
rect 20729 6273 20763 6307
rect 20821 6273 20855 6307
rect 20913 6273 20947 6307
rect 21070 6273 21104 6307
rect 21189 6273 21223 6307
rect 22477 6273 22511 6307
rect 8861 6205 8895 6239
rect 12449 6205 12483 6239
rect 13185 6205 13219 6239
rect 17141 6205 17175 6239
rect 17509 6205 17543 6239
rect 17969 6205 18003 6239
rect 15209 6137 15243 6171
rect 19901 6137 19935 6171
rect 12265 6069 12299 6103
rect 15025 6069 15059 6103
rect 16313 6069 16347 6103
rect 18153 6069 18187 6103
rect 20545 6069 20579 6103
rect 22201 6069 22235 6103
rect 12909 5865 12943 5899
rect 13093 5865 13127 5899
rect 16037 5865 16071 5899
rect 17141 5865 17175 5899
rect 17509 5865 17543 5899
rect 20729 5865 20763 5899
rect 21281 5865 21315 5899
rect 21649 5865 21683 5899
rect 22477 5865 22511 5899
rect 20545 5797 20579 5831
rect 16221 5729 16255 5763
rect 16313 5729 16347 5763
rect 20269 5729 20303 5763
rect 21465 5729 21499 5763
rect 13369 5661 13403 5695
rect 16681 5661 16715 5695
rect 17601 5661 17635 5695
rect 21189 5661 21223 5695
rect 21557 5661 21591 5695
rect 22569 5661 22603 5695
rect 16497 5525 16531 5559
rect 16589 5525 16623 5559
rect 22109 5525 22143 5559
rect 17049 5321 17083 5355
rect 20637 5321 20671 5355
rect 21281 5321 21315 5355
rect 21189 5253 21223 5287
rect 16865 5185 16899 5219
rect 17049 5185 17083 5219
rect 20177 5185 20211 5219
rect 21097 5185 21131 5219
rect 21373 5185 21407 5219
rect 20269 4981 20303 5015
<< metal1 >>
rect 5350 20816 5356 20868
rect 5408 20856 5414 20868
rect 10134 20856 10140 20868
rect 5408 20828 10140 20856
rect 5408 20816 5414 20828
rect 10134 20816 10140 20828
rect 10192 20816 10198 20868
rect 4890 20748 4896 20800
rect 4948 20788 4954 20800
rect 15838 20788 15844 20800
rect 4948 20760 15844 20788
rect 4948 20748 4954 20760
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 1104 20698 32632 20720
rect 1104 20646 8792 20698
rect 8844 20646 8856 20698
rect 8908 20646 8920 20698
rect 8972 20646 8984 20698
rect 9036 20646 9048 20698
rect 9100 20646 16634 20698
rect 16686 20646 16698 20698
rect 16750 20646 16762 20698
rect 16814 20646 16826 20698
rect 16878 20646 16890 20698
rect 16942 20646 24476 20698
rect 24528 20646 24540 20698
rect 24592 20646 24604 20698
rect 24656 20646 24668 20698
rect 24720 20646 24732 20698
rect 24784 20646 32318 20698
rect 32370 20646 32382 20698
rect 32434 20646 32446 20698
rect 32498 20646 32510 20698
rect 32562 20646 32574 20698
rect 32626 20646 32632 20698
rect 1104 20624 32632 20646
rect 2133 20587 2191 20593
rect 2133 20553 2145 20587
rect 2179 20584 2191 20587
rect 4430 20584 4436 20596
rect 2179 20556 4436 20584
rect 2179 20553 2191 20556
rect 2133 20547 2191 20553
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4890 20544 4896 20596
rect 4948 20544 4954 20596
rect 8110 20544 8116 20596
rect 8168 20544 8174 20596
rect 9490 20544 9496 20596
rect 9548 20544 9554 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 13538 20544 13544 20596
rect 13596 20544 13602 20596
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 17034 20544 17040 20596
rect 17092 20544 17098 20596
rect 27157 20587 27215 20593
rect 27157 20584 27169 20587
rect 17144 20556 27169 20584
rect 2777 20519 2835 20525
rect 2777 20485 2789 20519
rect 2823 20516 2835 20519
rect 4798 20516 4804 20528
rect 2823 20488 4804 20516
rect 2823 20485 2835 20488
rect 2777 20479 2835 20485
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 7469 20519 7527 20525
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 9692 20516 9720 20544
rect 7515 20488 9720 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 11698 20476 11704 20528
rect 11756 20476 11762 20528
rect 15378 20516 15384 20528
rect 11808 20488 15384 20516
rect 3421 20451 3479 20457
rect 3421 20417 3433 20451
rect 3467 20448 3479 20451
rect 3467 20420 4660 20448
rect 3467 20417 3479 20420
rect 3421 20411 3479 20417
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20349 4307 20383
rect 4632 20380 4660 20420
rect 4706 20408 4712 20460
rect 4764 20408 4770 20460
rect 5810 20408 5816 20460
rect 5868 20408 5874 20460
rect 5994 20408 6000 20460
rect 6052 20408 6058 20460
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20417 7619 20451
rect 7561 20411 7619 20417
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 5534 20380 5540 20392
rect 4632 20352 5540 20380
rect 4249 20343 4307 20349
rect 4264 20312 4292 20343
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 6086 20312 6092 20324
rect 4264 20284 6092 20312
rect 6086 20272 6092 20284
rect 6144 20272 6150 20324
rect 6733 20315 6791 20321
rect 6733 20281 6745 20315
rect 6779 20312 6791 20315
rect 7576 20312 7604 20411
rect 8312 20380 8340 20411
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 10042 20408 10048 20460
rect 10100 20448 10106 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10100 20420 10425 20448
rect 10100 20408 10106 20420
rect 10413 20417 10425 20420
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 8312 20352 10088 20380
rect 9950 20312 9956 20324
rect 6779 20284 7512 20312
rect 7576 20284 9956 20312
rect 6779 20281 6791 20284
rect 6733 20275 6791 20281
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 6822 20244 6828 20256
rect 5951 20216 6828 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7484 20244 7512 20284
rect 9950 20272 9956 20284
rect 10008 20272 10014 20324
rect 8110 20244 8116 20256
rect 7484 20216 8116 20244
rect 8110 20204 8116 20216
rect 8168 20204 8174 20256
rect 10060 20244 10088 20352
rect 10134 20340 10140 20392
rect 10192 20380 10198 20392
rect 10778 20380 10784 20392
rect 10192 20352 10784 20380
rect 10192 20340 10198 20352
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 10226 20272 10232 20324
rect 10284 20312 10290 20324
rect 10321 20315 10379 20321
rect 10321 20312 10333 20315
rect 10284 20284 10333 20312
rect 10284 20272 10290 20284
rect 10321 20281 10333 20284
rect 10367 20281 10379 20315
rect 10321 20275 10379 20281
rect 10413 20315 10471 20321
rect 10413 20281 10425 20315
rect 10459 20312 10471 20315
rect 10888 20312 10916 20411
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 11808 20448 11836 20488
rect 15378 20476 15384 20488
rect 15436 20476 15442 20528
rect 17144 20516 17172 20556
rect 27157 20553 27169 20556
rect 27203 20553 27215 20587
rect 27157 20547 27215 20553
rect 15488 20488 17172 20516
rect 11020 20420 11836 20448
rect 11020 20408 11026 20420
rect 11974 20408 11980 20460
rect 12032 20408 12038 20460
rect 12158 20408 12164 20460
rect 12216 20408 12222 20460
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13688 20420 13737 20448
rect 13688 20408 13694 20420
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 15197 20451 15255 20457
rect 15197 20417 15209 20451
rect 15243 20417 15255 20451
rect 15197 20411 15255 20417
rect 10459 20284 10916 20312
rect 11057 20315 11115 20321
rect 10459 20281 10471 20284
rect 10413 20275 10471 20281
rect 11057 20281 11069 20315
rect 11103 20312 11115 20315
rect 13814 20312 13820 20324
rect 11103 20284 13820 20312
rect 11103 20281 11115 20284
rect 11057 20275 11115 20281
rect 13814 20272 13820 20284
rect 13872 20272 13878 20324
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 10060 20216 14841 20244
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 15212 20244 15240 20411
rect 15289 20383 15347 20389
rect 15289 20349 15301 20383
rect 15335 20349 15347 20383
rect 15289 20343 15347 20349
rect 15304 20312 15332 20343
rect 15378 20340 15384 20392
rect 15436 20380 15442 20392
rect 15488 20389 15516 20488
rect 17402 20476 17408 20528
rect 17460 20516 17466 20528
rect 19429 20519 19487 20525
rect 19429 20516 19441 20519
rect 17460 20488 19441 20516
rect 17460 20476 17466 20488
rect 19429 20485 19441 20488
rect 19475 20485 19487 20519
rect 19429 20479 19487 20485
rect 19797 20519 19855 20525
rect 19797 20485 19809 20519
rect 19843 20516 19855 20519
rect 20441 20519 20499 20525
rect 20441 20516 20453 20519
rect 19843 20488 20453 20516
rect 19843 20485 19855 20488
rect 19797 20479 19855 20485
rect 20441 20485 20453 20488
rect 20487 20485 20499 20519
rect 20441 20479 20499 20485
rect 28077 20519 28135 20525
rect 28077 20485 28089 20519
rect 28123 20516 28135 20519
rect 29978 20519 30036 20525
rect 29978 20516 29990 20519
rect 28123 20488 29990 20516
rect 28123 20485 28135 20488
rect 28077 20479 28135 20485
rect 29978 20485 29990 20488
rect 30024 20485 30036 20519
rect 29978 20479 30036 20485
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 15436 20352 15485 20380
rect 15436 20340 15442 20352
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 16316 20380 16344 20411
rect 16390 20408 16396 20460
rect 16448 20448 16454 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16448 20420 16865 20448
rect 16448 20408 16454 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 18598 20408 18604 20460
rect 18656 20448 18662 20460
rect 18693 20451 18751 20457
rect 18693 20448 18705 20451
rect 18656 20420 18705 20448
rect 18656 20408 18662 20420
rect 18693 20417 18705 20420
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 18966 20448 18972 20460
rect 18923 20420 18972 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20162 20448 20168 20460
rect 19935 20420 20168 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20254 20408 20260 20460
rect 20312 20448 20318 20460
rect 20349 20451 20407 20457
rect 20349 20448 20361 20451
rect 20312 20420 20361 20448
rect 20312 20408 20318 20420
rect 20349 20417 20361 20420
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20898 20448 20904 20460
rect 20579 20420 20904 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20448 23351 20451
rect 23566 20448 23572 20460
rect 23339 20420 23572 20448
rect 23339 20417 23351 20420
rect 23293 20411 23351 20417
rect 23566 20408 23572 20420
rect 23624 20448 23630 20460
rect 25593 20451 25651 20457
rect 25593 20448 25605 20451
rect 23624 20420 25605 20448
rect 23624 20408 23630 20420
rect 25593 20417 25605 20420
rect 25639 20417 25651 20451
rect 25593 20411 25651 20417
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20448 25743 20451
rect 26234 20448 26240 20460
rect 25731 20420 26240 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27798 20408 27804 20460
rect 27856 20408 27862 20460
rect 30466 20408 30472 20460
rect 30524 20448 30530 20460
rect 31573 20451 31631 20457
rect 31573 20448 31585 20451
rect 30524 20420 31585 20448
rect 30524 20408 30530 20420
rect 31573 20417 31585 20420
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 17494 20380 17500 20392
rect 16316 20352 17500 20380
rect 15473 20343 15531 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20349 19579 20383
rect 19521 20343 19579 20349
rect 17402 20312 17408 20324
rect 15304 20284 17408 20312
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 19536 20312 19564 20343
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 23201 20383 23259 20389
rect 23201 20380 23213 20383
rect 22152 20352 23213 20380
rect 22152 20340 22158 20352
rect 23201 20349 23213 20352
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 26016 20352 26065 20380
rect 26016 20340 26022 20352
rect 26053 20349 26065 20352
rect 26099 20349 26111 20383
rect 26053 20343 26111 20349
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20380 28687 20383
rect 28675 20352 29684 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 17696 20284 19564 20312
rect 15746 20244 15752 20256
rect 15212 20216 15752 20244
rect 14829 20207 14887 20213
rect 15746 20204 15752 20216
rect 15804 20244 15810 20256
rect 17696 20244 17724 20284
rect 23014 20272 23020 20324
rect 23072 20312 23078 20324
rect 25869 20315 25927 20321
rect 25869 20312 25881 20315
rect 23072 20284 25881 20312
rect 23072 20272 23078 20284
rect 25869 20281 25881 20284
rect 25915 20281 25927 20315
rect 25869 20275 25927 20281
rect 15804 20216 17724 20244
rect 18785 20247 18843 20253
rect 15804 20204 15810 20216
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 18874 20244 18880 20256
rect 18831 20216 18880 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 19613 20247 19671 20253
rect 19613 20213 19625 20247
rect 19659 20244 19671 20247
rect 20438 20244 20444 20256
rect 19659 20216 20444 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 23661 20247 23719 20253
rect 23661 20213 23673 20247
rect 23707 20244 23719 20247
rect 24946 20244 24952 20256
rect 23707 20216 24952 20244
rect 23707 20213 23719 20216
rect 23661 20207 23719 20213
rect 24946 20204 24952 20216
rect 25004 20204 25010 20256
rect 29178 20204 29184 20256
rect 29236 20204 29242 20256
rect 29656 20244 29684 20352
rect 29730 20340 29736 20392
rect 29788 20340 29794 20392
rect 31113 20247 31171 20253
rect 31113 20244 31125 20247
rect 29656 20216 31125 20244
rect 31113 20213 31125 20216
rect 31159 20213 31171 20247
rect 31113 20207 31171 20213
rect 31662 20204 31668 20256
rect 31720 20204 31726 20256
rect 1104 20154 32476 20176
rect 1104 20102 4871 20154
rect 4923 20102 4935 20154
rect 4987 20102 4999 20154
rect 5051 20102 5063 20154
rect 5115 20102 5127 20154
rect 5179 20102 12713 20154
rect 12765 20102 12777 20154
rect 12829 20102 12841 20154
rect 12893 20102 12905 20154
rect 12957 20102 12969 20154
rect 13021 20102 20555 20154
rect 20607 20102 20619 20154
rect 20671 20102 20683 20154
rect 20735 20102 20747 20154
rect 20799 20102 20811 20154
rect 20863 20102 28397 20154
rect 28449 20102 28461 20154
rect 28513 20102 28525 20154
rect 28577 20102 28589 20154
rect 28641 20102 28653 20154
rect 28705 20102 32476 20154
rect 1104 20080 32476 20102
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 4706 20040 4712 20052
rect 3467 20012 4712 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 4706 20000 4712 20012
rect 4764 20000 4770 20052
rect 5350 20000 5356 20052
rect 5408 20000 5414 20052
rect 5994 20000 6000 20052
rect 6052 20040 6058 20052
rect 6052 20012 8064 20040
rect 6052 20000 6058 20012
rect 8036 19972 8064 20012
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 13541 20043 13599 20049
rect 8260 20012 12434 20040
rect 8260 20000 8266 20012
rect 8570 19972 8576 19984
rect 8036 19944 8576 19972
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 12406 19972 12434 20012
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 14182 20040 14188 20052
rect 13587 20012 14188 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 15010 20040 15016 20052
rect 14936 20012 15016 20040
rect 14936 19981 14964 20012
rect 15010 20000 15016 20012
rect 15068 20040 15074 20052
rect 15068 20012 18368 20040
rect 15068 20000 15074 20012
rect 14553 19975 14611 19981
rect 14553 19972 14565 19975
rect 12406 19944 14565 19972
rect 14553 19941 14565 19944
rect 14599 19941 14611 19975
rect 14553 19935 14611 19941
rect 14921 19975 14979 19981
rect 14921 19941 14933 19975
rect 14967 19941 14979 19975
rect 14921 19935 14979 19941
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19904 2191 19907
rect 2958 19904 2964 19916
rect 2179 19876 2964 19904
rect 2179 19873 2191 19876
rect 2133 19867 2191 19873
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 15286 19904 15292 19916
rect 8260 19876 9260 19904
rect 8260 19864 8266 19876
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19836 2651 19839
rect 2639 19808 2774 19836
rect 2639 19805 2651 19808
rect 2593 19799 2651 19805
rect 2746 19768 2774 19808
rect 3234 19796 3240 19848
rect 3292 19796 3298 19848
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19836 4031 19839
rect 4062 19836 4068 19848
rect 4019 19808 4068 19836
rect 4019 19805 4031 19808
rect 3973 19799 4031 19805
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19836 5963 19839
rect 7006 19836 7012 19848
rect 5951 19808 7012 19836
rect 5951 19805 5963 19808
rect 5905 19799 5963 19805
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 8110 19836 8116 19848
rect 7147 19808 8116 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 8110 19796 8116 19808
rect 8168 19836 8174 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 8168 19808 9137 19836
rect 8168 19796 8174 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9232 19836 9260 19876
rect 10152 19876 15292 19904
rect 9381 19839 9439 19845
rect 9381 19836 9393 19839
rect 9232 19808 9393 19836
rect 9125 19799 9183 19805
rect 9381 19805 9393 19808
rect 9427 19805 9439 19839
rect 10152 19836 10180 19876
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 18340 19904 18368 20012
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19981 20043 20039 20049
rect 19981 20040 19993 20043
rect 19024 20012 19993 20040
rect 19024 20000 19030 20012
rect 19981 20009 19993 20012
rect 20027 20009 20039 20043
rect 19981 20003 20039 20009
rect 19996 19972 20024 20003
rect 20162 20000 20168 20052
rect 20220 20000 20226 20052
rect 20438 20000 20444 20052
rect 20496 20040 20502 20052
rect 20625 20043 20683 20049
rect 20625 20040 20637 20043
rect 20496 20012 20637 20040
rect 20496 20000 20502 20012
rect 20625 20009 20637 20012
rect 20671 20009 20683 20043
rect 20625 20003 20683 20009
rect 22094 20000 22100 20052
rect 22152 20000 22158 20052
rect 25869 20043 25927 20049
rect 25869 20009 25881 20043
rect 25915 20040 25927 20043
rect 27798 20040 27804 20052
rect 25915 20012 27804 20040
rect 25915 20009 25927 20012
rect 25869 20003 25927 20009
rect 27798 20000 27804 20012
rect 27856 20000 27862 20052
rect 20990 19972 20996 19984
rect 19996 19944 20996 19972
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 24581 19975 24639 19981
rect 24581 19972 24593 19975
rect 21100 19944 24593 19972
rect 18340 19876 20852 19904
rect 9381 19799 9439 19805
rect 9508 19808 10180 19836
rect 11057 19839 11115 19845
rect 2746 19740 3464 19768
rect 2774 19660 2780 19712
rect 2832 19660 2838 19712
rect 3436 19700 3464 19740
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 4218 19771 4276 19777
rect 4218 19768 4230 19771
rect 3568 19740 4230 19768
rect 3568 19728 3574 19740
rect 4218 19737 4230 19740
rect 4264 19737 4276 19771
rect 7346 19771 7404 19777
rect 7346 19768 7358 19771
rect 4218 19731 4276 19737
rect 6104 19740 7358 19768
rect 4338 19700 4344 19712
rect 3436 19672 4344 19700
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 6104 19709 6132 19740
rect 7346 19737 7358 19740
rect 7392 19737 7404 19771
rect 7346 19731 7404 19737
rect 8202 19728 8208 19780
rect 8260 19768 8266 19780
rect 9508 19768 9536 19808
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 11238 19836 11244 19848
rect 11103 19808 11244 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19836 11759 19839
rect 12158 19836 12164 19848
rect 11747 19808 12164 19836
rect 11747 19805 11759 19808
rect 11701 19799 11759 19805
rect 8260 19740 9536 19768
rect 8260 19728 8266 19740
rect 9674 19728 9680 19780
rect 9732 19768 9738 19780
rect 11716 19768 11744 19799
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 12618 19836 12624 19848
rect 12299 19808 12624 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 13722 19796 13728 19848
rect 13780 19796 13786 19848
rect 14734 19796 14740 19848
rect 14792 19796 14798 19848
rect 15013 19839 15071 19845
rect 15013 19805 15025 19839
rect 15059 19836 15071 19839
rect 15378 19836 15384 19848
rect 15059 19808 15384 19836
rect 15059 19805 15071 19808
rect 15013 19799 15071 19805
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19836 15531 19839
rect 17313 19839 17371 19845
rect 17313 19836 17325 19839
rect 15519 19808 17325 19836
rect 15519 19805 15531 19808
rect 15473 19799 15531 19805
rect 17313 19805 17325 19808
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 9732 19740 11744 19768
rect 9732 19728 9738 19740
rect 12066 19728 12072 19780
rect 12124 19768 12130 19780
rect 12124 19740 14596 19768
rect 12124 19728 12130 19740
rect 6089 19703 6147 19709
rect 6089 19669 6101 19703
rect 6135 19669 6147 19703
rect 6089 19663 6147 19669
rect 8478 19660 8484 19712
rect 8536 19700 8542 19712
rect 9306 19700 9312 19712
rect 8536 19672 9312 19700
rect 8536 19660 8542 19672
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 9582 19660 9588 19712
rect 9640 19700 9646 19712
rect 10505 19703 10563 19709
rect 10505 19700 10517 19703
rect 9640 19672 10517 19700
rect 9640 19660 9646 19672
rect 10505 19669 10517 19672
rect 10551 19700 10563 19703
rect 10962 19700 10968 19712
rect 10551 19672 10968 19700
rect 10551 19669 10563 19672
rect 10505 19663 10563 19669
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11146 19660 11152 19712
rect 11204 19660 11210 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 13538 19700 13544 19712
rect 11848 19672 13544 19700
rect 11848 19660 11854 19672
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 14568 19700 14596 19740
rect 14642 19728 14648 19780
rect 14700 19768 14706 19780
rect 15488 19768 15516 19799
rect 17402 19796 17408 19848
rect 17460 19836 17466 19848
rect 17569 19839 17627 19845
rect 17569 19836 17581 19839
rect 17460 19808 17581 19836
rect 17460 19796 17466 19808
rect 17569 19805 17581 19808
rect 17615 19805 17627 19839
rect 17569 19799 17627 19805
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 18748 19808 19533 19836
rect 18748 19796 18754 19808
rect 19521 19805 19533 19808
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 19794 19836 19800 19848
rect 19659 19808 19800 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 19978 19845 19984 19848
rect 19971 19839 19984 19845
rect 19971 19805 19983 19839
rect 20036 19836 20042 19848
rect 20824 19845 20852 19876
rect 21100 19845 21128 19944
rect 24581 19941 24593 19944
rect 24627 19941 24639 19975
rect 29454 19972 29460 19984
rect 24581 19935 24639 19941
rect 25700 19944 29460 19972
rect 22370 19864 22376 19916
rect 22428 19904 22434 19916
rect 22925 19907 22983 19913
rect 22925 19904 22937 19907
rect 22428 19876 22937 19904
rect 22428 19864 22434 19876
rect 22925 19873 22937 19876
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 24854 19864 24860 19916
rect 24912 19864 24918 19916
rect 20809 19839 20867 19845
rect 20036 19808 20071 19836
rect 19971 19799 19984 19805
rect 19978 19796 19984 19799
rect 20036 19796 20042 19808
rect 20809 19805 20821 19839
rect 20855 19805 20867 19839
rect 20809 19799 20867 19805
rect 21085 19839 21143 19845
rect 21085 19805 21097 19839
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 15746 19777 15752 19780
rect 15740 19768 15752 19777
rect 14700 19740 15516 19768
rect 15707 19740 15752 19768
rect 14700 19728 14706 19740
rect 15740 19731 15752 19740
rect 15746 19728 15752 19731
rect 15804 19728 15810 19780
rect 18598 19768 18604 19780
rect 16776 19740 18604 19768
rect 16776 19700 16804 19740
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 20070 19728 20076 19780
rect 20128 19768 20134 19780
rect 21100 19768 21128 19799
rect 22002 19796 22008 19848
rect 22060 19796 22066 19848
rect 22189 19839 22247 19845
rect 22189 19805 22201 19839
rect 22235 19836 22247 19839
rect 22278 19836 22284 19848
rect 22235 19808 22284 19836
rect 22235 19805 22247 19808
rect 22189 19799 22247 19805
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 23014 19796 23020 19848
rect 23072 19796 23078 19848
rect 24946 19796 24952 19848
rect 25004 19796 25010 19848
rect 25700 19845 25728 19944
rect 29454 19932 29460 19944
rect 29512 19932 29518 19984
rect 26786 19864 26792 19916
rect 26844 19864 26850 19916
rect 25685 19839 25743 19845
rect 25685 19805 25697 19839
rect 25731 19805 25743 19839
rect 25685 19799 25743 19805
rect 26694 19796 26700 19848
rect 26752 19796 26758 19848
rect 28074 19796 28080 19848
rect 28132 19796 28138 19848
rect 28350 19796 28356 19848
rect 28408 19836 28414 19848
rect 28537 19839 28595 19845
rect 28537 19836 28549 19839
rect 28408 19808 28549 19836
rect 28408 19796 28414 19808
rect 28537 19805 28549 19808
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30282 19836 30288 19848
rect 29788 19808 30288 19836
rect 29788 19796 29794 19808
rect 30282 19796 30288 19808
rect 30340 19796 30346 19848
rect 30926 19796 30932 19848
rect 30984 19836 30990 19848
rect 31573 19839 31631 19845
rect 31573 19836 31585 19839
rect 30984 19808 31585 19836
rect 30984 19796 30990 19808
rect 31573 19805 31585 19808
rect 31619 19805 31631 19839
rect 31573 19799 31631 19805
rect 31849 19839 31907 19845
rect 31849 19805 31861 19839
rect 31895 19836 31907 19839
rect 31938 19836 31944 19848
rect 31895 19808 31944 19836
rect 31895 19805 31907 19808
rect 31849 19799 31907 19805
rect 31938 19796 31944 19808
rect 31996 19796 32002 19848
rect 20128 19740 21128 19768
rect 29181 19771 29239 19777
rect 20128 19728 20134 19740
rect 29181 19737 29193 19771
rect 29227 19768 29239 19771
rect 29978 19771 30036 19777
rect 29978 19768 29990 19771
rect 29227 19740 29990 19768
rect 29227 19737 29239 19740
rect 29181 19731 29239 19737
rect 29978 19737 29990 19740
rect 30024 19737 30036 19771
rect 29978 19731 30036 19737
rect 14568 19672 16804 19700
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19700 16911 19703
rect 17034 19700 17040 19712
rect 16899 19672 17040 19700
rect 16899 19669 16911 19672
rect 16853 19663 16911 19669
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 18693 19703 18751 19709
rect 18693 19669 18705 19703
rect 18739 19700 18751 19703
rect 18782 19700 18788 19712
rect 18739 19672 18788 19700
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20898 19700 20904 19712
rect 20036 19672 20904 19700
rect 20036 19660 20042 19672
rect 20898 19660 20904 19672
rect 20956 19700 20962 19712
rect 20993 19703 21051 19709
rect 20993 19700 21005 19703
rect 20956 19672 21005 19700
rect 20956 19660 20962 19672
rect 20993 19669 21005 19672
rect 21039 19700 21051 19703
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 21039 19672 22661 19700
rect 21039 19669 21051 19672
rect 20993 19663 21051 19669
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 22649 19663 22707 19669
rect 25958 19660 25964 19712
rect 26016 19700 26022 19712
rect 26329 19703 26387 19709
rect 26329 19700 26341 19703
rect 26016 19672 26341 19700
rect 26016 19660 26022 19672
rect 26329 19669 26341 19672
rect 26375 19669 26387 19703
rect 26329 19663 26387 19669
rect 27890 19660 27896 19712
rect 27948 19660 27954 19712
rect 31113 19703 31171 19709
rect 31113 19669 31125 19703
rect 31159 19700 31171 19703
rect 31570 19700 31576 19712
rect 31159 19672 31576 19700
rect 31159 19669 31171 19672
rect 31113 19663 31171 19669
rect 31570 19660 31576 19672
rect 31628 19660 31634 19712
rect 1104 19610 32632 19632
rect 1104 19558 8792 19610
rect 8844 19558 8856 19610
rect 8908 19558 8920 19610
rect 8972 19558 8984 19610
rect 9036 19558 9048 19610
rect 9100 19558 16634 19610
rect 16686 19558 16698 19610
rect 16750 19558 16762 19610
rect 16814 19558 16826 19610
rect 16878 19558 16890 19610
rect 16942 19558 24476 19610
rect 24528 19558 24540 19610
rect 24592 19558 24604 19610
rect 24656 19558 24668 19610
rect 24720 19558 24732 19610
rect 24784 19558 32318 19610
rect 32370 19558 32382 19610
rect 32434 19558 32446 19610
rect 32498 19558 32510 19610
rect 32562 19558 32574 19610
rect 32626 19558 32632 19610
rect 1104 19536 32632 19558
rect 1762 19456 1768 19508
rect 1820 19456 1826 19508
rect 2409 19499 2467 19505
rect 2409 19465 2421 19499
rect 2455 19496 2467 19499
rect 3510 19496 3516 19508
rect 2455 19468 3516 19496
rect 2455 19465 2467 19468
rect 2409 19459 2467 19465
rect 3510 19456 3516 19468
rect 3568 19456 3574 19508
rect 6546 19456 6552 19508
rect 6604 19496 6610 19508
rect 9125 19499 9183 19505
rect 9125 19496 9137 19499
rect 6604 19468 9137 19496
rect 6604 19456 6610 19468
rect 9125 19465 9137 19468
rect 9171 19465 9183 19499
rect 9125 19459 9183 19465
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 9732 19468 10517 19496
rect 9732 19456 9738 19468
rect 10505 19465 10517 19468
rect 10551 19465 10563 19499
rect 10505 19459 10563 19465
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 16025 19499 16083 19505
rect 12216 19468 12848 19496
rect 12216 19456 12222 19468
rect 2774 19388 2780 19440
rect 2832 19428 2838 19440
rect 4402 19431 4460 19437
rect 4402 19428 4414 19431
rect 2832 19400 4414 19428
rect 2832 19388 2838 19400
rect 4402 19397 4414 19400
rect 4448 19397 4460 19431
rect 7837 19431 7895 19437
rect 7837 19428 7849 19431
rect 4402 19391 4460 19397
rect 6840 19400 7849 19428
rect 6840 19372 6868 19400
rect 7837 19397 7849 19400
rect 7883 19428 7895 19431
rect 9030 19428 9036 19440
rect 7883 19400 9036 19428
rect 7883 19397 7895 19400
rect 7837 19391 7895 19397
rect 9030 19388 9036 19400
rect 9088 19388 9094 19440
rect 9214 19388 9220 19440
rect 9272 19437 9278 19440
rect 9272 19431 9335 19437
rect 9272 19397 9289 19431
rect 9323 19397 9335 19431
rect 9272 19391 9335 19397
rect 9272 19388 9278 19391
rect 9490 19388 9496 19440
rect 9548 19388 9554 19440
rect 10042 19388 10048 19440
rect 10100 19428 10106 19440
rect 10100 19400 10916 19428
rect 10100 19388 10106 19400
rect 10888 19372 10916 19400
rect 11146 19388 11152 19440
rect 11204 19428 11210 19440
rect 11204 19400 12388 19428
rect 11204 19388 11210 19400
rect 2222 19320 2228 19372
rect 2280 19320 2286 19372
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19360 3111 19363
rect 3142 19360 3148 19372
rect 3099 19332 3148 19360
rect 3099 19329 3111 19332
rect 3053 19323 3111 19329
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3418 19360 3424 19372
rect 3375 19332 3424 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 2866 19252 2872 19304
rect 2924 19252 2930 19304
rect 2958 19252 2964 19304
rect 3016 19292 3022 19304
rect 3252 19292 3280 19323
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 6822 19320 6828 19372
rect 6880 19320 6886 19372
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 7098 19360 7104 19372
rect 7055 19332 7104 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7098 19320 7104 19332
rect 7156 19360 7162 19372
rect 7653 19363 7711 19369
rect 7653 19360 7665 19363
rect 7156 19332 7665 19360
rect 7156 19320 7162 19332
rect 7653 19329 7665 19332
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 3970 19292 3976 19304
rect 3016 19264 3976 19292
rect 3016 19252 3022 19264
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4154 19252 4160 19304
rect 4212 19252 4218 19304
rect 7668 19292 7696 19323
rect 8018 19320 8024 19372
rect 8076 19360 8082 19372
rect 8202 19360 8208 19372
rect 8076 19332 8208 19360
rect 8076 19320 8082 19332
rect 8202 19320 8208 19332
rect 8260 19360 8266 19372
rect 8297 19363 8355 19369
rect 8297 19360 8309 19363
rect 8260 19332 8309 19360
rect 8260 19320 8266 19332
rect 8297 19329 8309 19332
rect 8343 19329 8355 19363
rect 8297 19323 8355 19329
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 8570 19360 8576 19372
rect 8527 19332 8576 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 8570 19320 8576 19332
rect 8628 19360 8634 19372
rect 9582 19360 9588 19372
rect 8628 19332 9588 19360
rect 8628 19320 8634 19332
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 9950 19320 9956 19372
rect 10008 19360 10014 19372
rect 10410 19360 10416 19372
rect 10008 19332 10416 19360
rect 10008 19320 10014 19332
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 10870 19320 10876 19372
rect 10928 19320 10934 19372
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 12360 19369 12388 19400
rect 12820 19369 12848 19468
rect 16025 19465 16037 19499
rect 16071 19496 16083 19499
rect 16390 19496 16396 19508
rect 16071 19468 16396 19496
rect 16071 19465 16083 19468
rect 16025 19459 16083 19465
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 17037 19499 17095 19505
rect 17037 19465 17049 19499
rect 17083 19496 17095 19499
rect 17126 19496 17132 19508
rect 17083 19468 17132 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 18598 19456 18604 19508
rect 18656 19456 18662 19508
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19935 19468 20453 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20441 19465 20453 19468
rect 20487 19496 20499 19499
rect 20898 19496 20904 19508
rect 20487 19468 20904 19496
rect 20487 19465 20499 19468
rect 20441 19459 20499 19465
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 20990 19456 20996 19508
rect 21048 19496 21054 19508
rect 21361 19499 21419 19505
rect 21361 19496 21373 19499
rect 21048 19468 21373 19496
rect 21048 19456 21054 19468
rect 21361 19465 21373 19468
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 25409 19499 25467 19505
rect 25409 19465 25421 19499
rect 25455 19496 25467 19499
rect 26694 19496 26700 19508
rect 25455 19468 26700 19496
rect 25455 19465 25467 19468
rect 25409 19459 25467 19465
rect 26694 19456 26700 19468
rect 26752 19456 26758 19508
rect 26786 19456 26792 19508
rect 26844 19496 26850 19508
rect 27157 19499 27215 19505
rect 27157 19496 27169 19499
rect 26844 19468 27169 19496
rect 26844 19456 26850 19468
rect 27157 19465 27169 19468
rect 27203 19465 27215 19499
rect 27157 19459 27215 19465
rect 28350 19456 28356 19508
rect 28408 19456 28414 19508
rect 29178 19456 29184 19508
rect 29236 19496 29242 19508
rect 29236 19468 29868 19496
rect 29236 19456 29242 19468
rect 13078 19388 13084 19440
rect 13136 19428 13142 19440
rect 13817 19431 13875 19437
rect 13817 19428 13829 19431
rect 13136 19400 13829 19428
rect 13136 19388 13142 19400
rect 13817 19397 13829 19400
rect 13863 19397 13875 19431
rect 13817 19391 13875 19397
rect 15286 19388 15292 19440
rect 15344 19428 15350 19440
rect 22186 19428 22192 19440
rect 15344 19400 17908 19428
rect 15344 19388 15350 19400
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 12805 19363 12863 19369
rect 12805 19329 12817 19363
rect 12851 19329 12863 19363
rect 12805 19323 12863 19329
rect 13170 19320 13176 19372
rect 13228 19320 13234 19372
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 13541 19363 13599 19369
rect 13541 19360 13553 19363
rect 13504 19332 13553 19360
rect 13504 19320 13510 19332
rect 13541 19329 13553 19332
rect 13587 19329 13599 19363
rect 13541 19323 13599 19329
rect 14642 19320 14648 19372
rect 14700 19320 14706 19372
rect 14912 19363 14970 19369
rect 14912 19329 14924 19363
rect 14958 19360 14970 19363
rect 16482 19360 16488 19372
rect 14958 19332 16488 19360
rect 14958 19329 14970 19332
rect 14912 19323 14970 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 17034 19360 17040 19372
rect 16899 19332 17040 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17880 19369 17908 19400
rect 18064 19400 22192 19428
rect 18064 19369 18092 19400
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 18049 19363 18107 19369
rect 17911 19332 18000 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 17972 19292 18000 19332
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 18156 19332 18736 19360
rect 18156 19292 18184 19332
rect 7668 19264 14688 19292
rect 17972 19264 18184 19292
rect 18708 19292 18736 19332
rect 18782 19320 18788 19372
rect 18840 19320 18846 19372
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19360 19487 19363
rect 19518 19360 19524 19372
rect 19475 19332 19524 19360
rect 19475 19329 19487 19332
rect 19429 19323 19487 19329
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 20346 19320 20352 19372
rect 20404 19320 20410 19372
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 21468 19369 21496 19400
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 25866 19428 25872 19440
rect 25240 19400 25872 19428
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20496 19332 20637 19360
rect 20496 19320 20502 19332
rect 20625 19329 20637 19332
rect 20671 19329 20683 19363
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 20625 19323 20683 19329
rect 20732 19332 21281 19360
rect 20162 19292 20168 19304
rect 18708 19264 20168 19292
rect 5537 19227 5595 19233
rect 5537 19193 5549 19227
rect 5583 19224 5595 19227
rect 5810 19224 5816 19236
rect 5583 19196 5816 19224
rect 5583 19193 5595 19196
rect 5537 19187 5595 19193
rect 5810 19184 5816 19196
rect 5868 19224 5874 19236
rect 8018 19224 8024 19236
rect 5868 19196 8024 19224
rect 5868 19184 5874 19196
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 14458 19224 14464 19236
rect 9640 19196 14464 19224
rect 9640 19184 9646 19196
rect 14458 19184 14464 19196
rect 14516 19184 14522 19236
rect 6914 19116 6920 19168
rect 6972 19116 6978 19168
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 7469 19159 7527 19165
rect 7469 19156 7481 19159
rect 7248 19128 7481 19156
rect 7248 19116 7254 19128
rect 7469 19125 7481 19128
rect 7515 19125 7527 19159
rect 7469 19119 7527 19125
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 9030 19116 9036 19168
rect 9088 19156 9094 19168
rect 9309 19159 9367 19165
rect 9309 19156 9321 19159
rect 9088 19128 9321 19156
rect 9088 19116 9094 19128
rect 9309 19125 9321 19128
rect 9355 19125 9367 19159
rect 9309 19119 9367 19125
rect 9398 19116 9404 19168
rect 9456 19156 9462 19168
rect 14550 19156 14556 19168
rect 9456 19128 14556 19156
rect 9456 19116 9462 19128
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 14660 19156 14688 19264
rect 20162 19252 20168 19264
rect 20220 19292 20226 19304
rect 20732 19292 20760 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 22152 19332 22416 19360
rect 22152 19320 22158 19332
rect 20220 19264 20760 19292
rect 20220 19252 20226 19264
rect 21174 19252 21180 19304
rect 21232 19292 21238 19304
rect 22002 19292 22008 19304
rect 21232 19264 22008 19292
rect 21232 19252 21238 19264
rect 22002 19252 22008 19264
rect 22060 19292 22066 19304
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 22060 19264 22201 19292
rect 22060 19252 22066 19264
rect 22189 19261 22201 19264
rect 22235 19261 22247 19295
rect 22189 19255 22247 19261
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 22388 19301 22416 19332
rect 23198 19320 23204 19372
rect 23256 19320 23262 19372
rect 25240 19369 25268 19400
rect 25866 19388 25872 19400
rect 25924 19388 25930 19440
rect 27430 19428 27436 19440
rect 26344 19400 27436 19428
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 23584 19332 24225 19360
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19261 22431 19295
rect 22373 19255 22431 19261
rect 22465 19295 22523 19301
rect 22465 19261 22477 19295
rect 22511 19292 22523 19295
rect 22738 19292 22744 19304
rect 22511 19264 22744 19292
rect 22511 19261 22523 19264
rect 22465 19255 22523 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 17957 19227 18015 19233
rect 17957 19193 17969 19227
rect 18003 19224 18015 19227
rect 18690 19224 18696 19236
rect 18003 19196 18696 19224
rect 18003 19193 18015 19196
rect 17957 19187 18015 19193
rect 18690 19184 18696 19196
rect 18748 19184 18754 19236
rect 20809 19227 20867 19233
rect 20809 19193 20821 19227
rect 20855 19224 20867 19227
rect 23124 19224 23152 19255
rect 23584 19233 23612 19332
rect 24213 19329 24225 19332
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 25409 19363 25467 19369
rect 25409 19329 25421 19363
rect 25455 19360 25467 19363
rect 26234 19360 26240 19372
rect 25455 19332 26240 19360
rect 25455 19329 25467 19332
rect 25409 19323 25467 19329
rect 26234 19320 26240 19332
rect 26292 19320 26298 19372
rect 26344 19369 26372 19400
rect 27430 19388 27436 19400
rect 27488 19388 27494 19440
rect 28810 19388 28816 19440
rect 28868 19428 28874 19440
rect 29840 19428 29868 19468
rect 31478 19456 31484 19508
rect 31536 19496 31542 19508
rect 31665 19499 31723 19505
rect 31665 19496 31677 19499
rect 31536 19468 31677 19496
rect 31536 19456 31542 19468
rect 31665 19465 31677 19468
rect 31711 19465 31723 19499
rect 31665 19459 31723 19465
rect 30530 19431 30588 19437
rect 30530 19428 30542 19431
rect 28868 19400 29776 19428
rect 29840 19400 30542 19428
rect 28868 19388 28874 19400
rect 26329 19363 26387 19369
rect 26329 19329 26341 19363
rect 26375 19329 26387 19363
rect 26329 19323 26387 19329
rect 26510 19320 26516 19372
rect 26568 19360 26574 19372
rect 27525 19363 27583 19369
rect 27525 19360 27537 19363
rect 26568 19332 27537 19360
rect 26568 19320 26574 19332
rect 27525 19329 27537 19332
rect 27571 19329 27583 19363
rect 27525 19323 27583 19329
rect 27890 19320 27896 19372
rect 27948 19360 27954 19372
rect 29748 19369 29776 19400
rect 30530 19397 30542 19400
rect 30576 19397 30588 19431
rect 30530 19391 30588 19397
rect 29466 19363 29524 19369
rect 29466 19360 29478 19363
rect 27948 19332 29478 19360
rect 27948 19320 27954 19332
rect 29466 19329 29478 19332
rect 29512 19329 29524 19363
rect 29466 19323 29524 19329
rect 29733 19363 29791 19369
rect 29733 19329 29745 19363
rect 29779 19360 29791 19363
rect 30285 19363 30343 19369
rect 30285 19360 30297 19363
rect 29779 19332 30297 19360
rect 29779 19329 29791 19332
rect 29733 19323 29791 19329
rect 30285 19329 30297 19332
rect 30331 19329 30343 19363
rect 30285 19323 30343 19329
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 25958 19292 25964 19304
rect 24351 19264 25964 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 25958 19252 25964 19264
rect 26016 19252 26022 19304
rect 26418 19252 26424 19304
rect 26476 19292 26482 19304
rect 27433 19295 27491 19301
rect 27433 19292 27445 19295
rect 26476 19264 27445 19292
rect 26476 19252 26482 19264
rect 27433 19261 27445 19264
rect 27479 19261 27491 19295
rect 27433 19255 27491 19261
rect 20855 19196 23152 19224
rect 23569 19227 23627 19233
rect 20855 19193 20867 19196
rect 20809 19187 20867 19193
rect 23569 19193 23581 19227
rect 23615 19193 23627 19227
rect 23569 19187 23627 19193
rect 24581 19227 24639 19233
rect 24581 19193 24593 19227
rect 24627 19224 24639 19227
rect 24854 19224 24860 19236
rect 24627 19196 24860 19224
rect 24627 19193 24639 19196
rect 24581 19187 24639 19193
rect 24854 19184 24860 19196
rect 24912 19184 24918 19236
rect 25866 19184 25872 19236
rect 25924 19184 25930 19236
rect 15838 19156 15844 19168
rect 14660 19128 15844 19156
rect 15838 19116 15844 19128
rect 15896 19156 15902 19168
rect 17126 19156 17132 19168
rect 15896 19128 17132 19156
rect 15896 19116 15902 19128
rect 17126 19116 17132 19128
rect 17184 19116 17190 19168
rect 18414 19116 18420 19168
rect 18472 19156 18478 19168
rect 19521 19159 19579 19165
rect 19521 19156 19533 19159
rect 18472 19128 19533 19156
rect 18472 19116 18478 19128
rect 19521 19125 19533 19128
rect 19567 19156 19579 19159
rect 19702 19156 19708 19168
rect 19567 19128 19708 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 22002 19116 22008 19168
rect 22060 19116 22066 19168
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 26053 19159 26111 19165
rect 26053 19156 26065 19159
rect 22704 19128 26065 19156
rect 22704 19116 22710 19128
rect 26053 19125 26065 19128
rect 26099 19156 26111 19159
rect 26326 19156 26332 19168
rect 26099 19128 26332 19156
rect 26099 19125 26111 19128
rect 26053 19119 26111 19125
rect 26326 19116 26332 19128
rect 26384 19156 26390 19168
rect 27338 19156 27344 19168
rect 26384 19128 27344 19156
rect 26384 19116 26390 19128
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 1104 19066 32476 19088
rect 1104 19014 4871 19066
rect 4923 19014 4935 19066
rect 4987 19014 4999 19066
rect 5051 19014 5063 19066
rect 5115 19014 5127 19066
rect 5179 19014 12713 19066
rect 12765 19014 12777 19066
rect 12829 19014 12841 19066
rect 12893 19014 12905 19066
rect 12957 19014 12969 19066
rect 13021 19014 20555 19066
rect 20607 19014 20619 19066
rect 20671 19014 20683 19066
rect 20735 19014 20747 19066
rect 20799 19014 20811 19066
rect 20863 19014 28397 19066
rect 28449 19014 28461 19066
rect 28513 19014 28525 19066
rect 28577 19014 28589 19066
rect 28641 19014 28653 19066
rect 28705 19014 32476 19066
rect 1104 18992 32476 19014
rect 2590 18912 2596 18964
rect 2648 18952 2654 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2648 18924 2973 18952
rect 2648 18912 2654 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 2961 18915 3019 18921
rect 4157 18955 4215 18961
rect 4157 18921 4169 18955
rect 4203 18952 4215 18955
rect 4338 18952 4344 18964
rect 4203 18924 4344 18952
rect 4203 18921 4215 18924
rect 4157 18915 4215 18921
rect 4338 18912 4344 18924
rect 4396 18912 4402 18964
rect 5537 18955 5595 18961
rect 5537 18921 5549 18955
rect 5583 18952 5595 18955
rect 7098 18952 7104 18964
rect 5583 18924 7104 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 8478 18952 8484 18964
rect 7208 18924 8484 18952
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 2777 18887 2835 18893
rect 2777 18884 2789 18887
rect 2280 18856 2789 18884
rect 2280 18844 2286 18856
rect 2777 18853 2789 18856
rect 2823 18853 2835 18887
rect 2777 18847 2835 18853
rect 4062 18844 4068 18896
rect 4120 18884 4126 18896
rect 4249 18887 4307 18893
rect 4249 18884 4261 18887
rect 4120 18856 4261 18884
rect 4120 18844 4126 18856
rect 4249 18853 4261 18856
rect 4295 18853 4307 18887
rect 4249 18847 4307 18853
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 5810 18816 5816 18828
rect 4663 18788 5816 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 7208 18816 7236 18924
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 8662 18912 8668 18964
rect 8720 18952 8726 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8720 18924 9229 18952
rect 8720 18912 8726 18924
rect 9217 18921 9229 18924
rect 9263 18952 9275 18955
rect 9490 18952 9496 18964
rect 9263 18924 9496 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 10928 18924 12296 18952
rect 10928 18912 10934 18924
rect 11054 18844 11060 18896
rect 11112 18884 11118 18896
rect 11701 18887 11759 18893
rect 11701 18884 11713 18887
rect 11112 18856 11713 18884
rect 11112 18844 11118 18856
rect 11701 18853 11713 18856
rect 11747 18884 11759 18887
rect 11882 18884 11888 18896
rect 11747 18856 11888 18884
rect 11747 18853 11759 18856
rect 11701 18847 11759 18853
rect 11882 18844 11888 18856
rect 11940 18844 11946 18896
rect 6012 18788 7236 18816
rect 2130 18708 2136 18760
rect 2188 18708 2194 18760
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 2958 18748 2964 18760
rect 2363 18720 2964 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 3329 18751 3387 18757
rect 3329 18717 3341 18751
rect 3375 18748 3387 18751
rect 3418 18748 3424 18760
rect 3375 18720 3424 18748
rect 3375 18717 3387 18720
rect 3329 18711 3387 18717
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18748 5687 18751
rect 6012 18748 6040 18788
rect 10594 18776 10600 18828
rect 10652 18816 10658 18828
rect 12268 18816 12296 18924
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 17402 18952 17408 18964
rect 14608 18924 17408 18952
rect 14608 18912 14614 18924
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 18690 18912 18696 18964
rect 18748 18912 18754 18964
rect 18785 18955 18843 18961
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 20254 18952 20260 18964
rect 18831 18924 20260 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 20254 18912 20260 18924
rect 20312 18912 20318 18964
rect 21174 18912 21180 18964
rect 21232 18912 21238 18964
rect 21266 18912 21272 18964
rect 21324 18952 21330 18964
rect 21324 18924 26096 18952
rect 21324 18912 21330 18924
rect 13446 18844 13452 18896
rect 13504 18884 13510 18896
rect 17221 18887 17279 18893
rect 13504 18856 16804 18884
rect 13504 18844 13510 18856
rect 12437 18819 12495 18825
rect 12437 18816 12449 18819
rect 10652 18788 12204 18816
rect 12268 18788 12449 18816
rect 10652 18776 10658 18788
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 5675 18720 6040 18748
rect 6104 18720 6285 18748
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 2222 18572 2228 18624
rect 2280 18572 2286 18624
rect 2866 18572 2872 18624
rect 2924 18612 2930 18624
rect 2961 18615 3019 18621
rect 2961 18612 2973 18615
rect 2924 18584 2973 18612
rect 2924 18572 2930 18584
rect 2961 18581 2973 18584
rect 3007 18612 3019 18615
rect 4062 18612 4068 18624
rect 3007 18584 4068 18612
rect 3007 18581 3019 18584
rect 2961 18575 3019 18581
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 6104 18612 6132 18720
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 8168 18720 8217 18748
rect 8168 18708 8174 18720
rect 8205 18717 8217 18720
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8352 18720 9137 18748
rect 8352 18708 8358 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 6181 18683 6239 18689
rect 6181 18649 6193 18683
rect 6227 18680 6239 18683
rect 7960 18683 8018 18689
rect 6227 18652 7880 18680
rect 6227 18649 6239 18652
rect 6181 18643 6239 18649
rect 6825 18615 6883 18621
rect 6825 18612 6837 18615
rect 6104 18584 6837 18612
rect 6825 18581 6837 18584
rect 6871 18612 6883 18615
rect 7098 18612 7104 18624
rect 6871 18584 7104 18612
rect 6871 18581 6883 18584
rect 6825 18575 6883 18581
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 7852 18612 7880 18652
rect 7960 18649 7972 18683
rect 8006 18680 8018 18683
rect 8662 18680 8668 18692
rect 8006 18652 8668 18680
rect 8006 18649 8018 18652
rect 7960 18643 8018 18649
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 9140 18680 9168 18711
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 9490 18748 9496 18760
rect 9364 18720 9496 18748
rect 9364 18708 9370 18720
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18748 9643 18751
rect 9674 18748 9680 18760
rect 9631 18720 9680 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 10410 18708 10416 18760
rect 10468 18748 10474 18760
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 10468 18720 10977 18748
rect 10468 18708 10474 18720
rect 10965 18717 10977 18720
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 12176 18757 12204 18788
rect 12437 18785 12449 18788
rect 12483 18785 12495 18819
rect 12437 18779 12495 18785
rect 14734 18776 14740 18828
rect 14792 18816 14798 18828
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 14792 18788 14841 18816
rect 14792 18776 14798 18788
rect 14829 18785 14841 18788
rect 14875 18785 14887 18819
rect 14829 18779 14887 18785
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 16776 18816 16804 18856
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 19610 18884 19616 18896
rect 17267 18856 19616 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 19610 18844 19616 18856
rect 19668 18844 19674 18896
rect 19702 18844 19708 18896
rect 19760 18844 19766 18896
rect 19794 18844 19800 18896
rect 19852 18884 19858 18896
rect 19852 18856 21956 18884
rect 19852 18844 19858 18856
rect 15243 18788 16712 18816
rect 16776 18788 17356 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 11112 18720 11621 18748
rect 11112 18708 11118 18720
rect 11609 18717 11621 18720
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 10781 18683 10839 18689
rect 10781 18680 10793 18683
rect 9140 18652 10793 18680
rect 10781 18649 10793 18652
rect 10827 18649 10839 18683
rect 10781 18643 10839 18649
rect 9398 18612 9404 18624
rect 7852 18584 9404 18612
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 9769 18615 9827 18621
rect 9769 18581 9781 18615
rect 9815 18612 9827 18615
rect 9950 18612 9956 18624
rect 9815 18584 9956 18612
rect 9815 18581 9827 18584
rect 9769 18575 9827 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10796 18612 10824 18643
rect 11146 18640 11152 18692
rect 11204 18640 11210 18692
rect 11330 18612 11336 18624
rect 10796 18584 11336 18612
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 11624 18612 11652 18711
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 13262 18748 13268 18760
rect 12584 18720 13268 18748
rect 12584 18708 12590 18720
rect 13262 18708 13268 18720
rect 13320 18708 13326 18760
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 13078 18640 13084 18692
rect 13136 18680 13142 18692
rect 13464 18680 13492 18711
rect 13538 18708 13544 18760
rect 13596 18708 13602 18760
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 15657 18751 15715 18757
rect 15657 18748 15669 18751
rect 15528 18720 15669 18748
rect 15528 18708 15534 18720
rect 15657 18717 15669 18720
rect 15703 18717 15715 18751
rect 15657 18711 15715 18717
rect 15838 18708 15844 18760
rect 15896 18708 15902 18760
rect 15930 18708 15936 18760
rect 15988 18748 15994 18760
rect 16684 18757 16712 18788
rect 16669 18751 16727 18757
rect 15988 18720 16620 18748
rect 15988 18708 15994 18720
rect 13136 18652 13492 18680
rect 15028 18680 15056 18708
rect 15562 18680 15568 18692
rect 15028 18652 15568 18680
rect 13136 18640 13142 18652
rect 15562 18640 15568 18652
rect 15620 18640 15626 18692
rect 12434 18612 12440 18624
rect 11624 18584 12440 18612
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 13173 18615 13231 18621
rect 13173 18612 13185 18615
rect 12768 18584 13185 18612
rect 12768 18572 12774 18584
rect 13173 18581 13185 18584
rect 13219 18581 13231 18615
rect 13173 18575 13231 18581
rect 14458 18572 14464 18624
rect 14516 18612 14522 18624
rect 15838 18612 15844 18624
rect 14516 18584 15844 18612
rect 14516 18572 14522 18584
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16025 18615 16083 18621
rect 16025 18581 16037 18615
rect 16071 18612 16083 18615
rect 16298 18612 16304 18624
rect 16071 18584 16304 18612
rect 16071 18581 16083 18584
rect 16025 18575 16083 18581
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16482 18572 16488 18624
rect 16540 18572 16546 18624
rect 16592 18612 16620 18720
rect 16669 18717 16681 18751
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 17126 18708 17132 18760
rect 17184 18708 17190 18760
rect 17328 18757 17356 18788
rect 18874 18776 18880 18828
rect 18932 18776 18938 18828
rect 21928 18825 21956 18856
rect 22370 18844 22376 18896
rect 22428 18844 22434 18896
rect 23566 18844 23572 18896
rect 23624 18844 23630 18896
rect 26068 18825 26096 18924
rect 26510 18912 26516 18964
rect 26568 18912 26574 18964
rect 27341 18955 27399 18961
rect 27341 18921 27353 18955
rect 27387 18952 27399 18955
rect 27430 18952 27436 18964
rect 27387 18924 27436 18952
rect 27387 18921 27399 18924
rect 27341 18915 27399 18921
rect 27430 18912 27436 18924
rect 27488 18912 27494 18964
rect 28074 18912 28080 18964
rect 28132 18912 28138 18964
rect 28997 18955 29055 18961
rect 28997 18921 29009 18955
rect 29043 18952 29055 18955
rect 30466 18952 30472 18964
rect 29043 18924 30472 18952
rect 29043 18921 29055 18924
rect 28997 18915 29055 18921
rect 30466 18912 30472 18924
rect 30524 18912 30530 18964
rect 26234 18844 26240 18896
rect 26292 18884 26298 18896
rect 26973 18887 27031 18893
rect 26973 18884 26985 18887
rect 26292 18856 26985 18884
rect 26292 18844 26298 18856
rect 26973 18853 26985 18856
rect 27019 18853 27031 18887
rect 26973 18847 27031 18853
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18785 19947 18819
rect 19889 18779 19947 18785
rect 21913 18819 21971 18825
rect 21913 18785 21925 18819
rect 21959 18785 21971 18819
rect 21913 18779 21971 18785
rect 26053 18819 26111 18825
rect 26053 18785 26065 18819
rect 26099 18785 26111 18819
rect 26053 18779 26111 18785
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 18601 18751 18659 18757
rect 18601 18748 18613 18751
rect 18564 18720 18613 18748
rect 18564 18708 18570 18720
rect 18601 18717 18613 18720
rect 18647 18717 18659 18751
rect 19904 18748 19932 18779
rect 20438 18748 20444 18760
rect 19904 18720 20444 18748
rect 18601 18711 18659 18717
rect 20438 18708 20444 18720
rect 20496 18748 20502 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 20496 18720 20545 18748
rect 20496 18708 20502 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 20626 18751 20684 18757
rect 20626 18717 20638 18751
rect 20672 18717 20684 18751
rect 20626 18711 20684 18717
rect 19429 18683 19487 18689
rect 19429 18649 19441 18683
rect 19475 18680 19487 18683
rect 19518 18680 19524 18692
rect 19475 18652 19524 18680
rect 19475 18649 19487 18652
rect 19429 18643 19487 18649
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 20346 18640 20352 18692
rect 20404 18680 20410 18692
rect 20640 18680 20668 18711
rect 20806 18708 20812 18760
rect 20864 18708 20870 18760
rect 21039 18751 21097 18757
rect 21039 18748 21051 18751
rect 21013 18717 21051 18748
rect 21085 18748 21097 18751
rect 21266 18748 21272 18760
rect 21085 18720 21272 18748
rect 21085 18717 21097 18720
rect 21013 18711 21097 18717
rect 20404 18652 20668 18680
rect 20404 18640 20410 18652
rect 20898 18640 20904 18692
rect 20956 18640 20962 18692
rect 18874 18612 18880 18624
rect 16592 18584 18880 18612
rect 18874 18572 18880 18584
rect 18932 18612 18938 18624
rect 21013 18612 21041 18711
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 22002 18708 22008 18760
rect 22060 18708 22066 18760
rect 23198 18708 23204 18760
rect 23256 18748 23262 18760
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 23256 18720 23305 18748
rect 23256 18708 23262 18720
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 24394 18748 24400 18760
rect 23293 18711 23351 18717
rect 23492 18720 24400 18748
rect 21450 18640 21456 18692
rect 21508 18680 21514 18692
rect 23492 18680 23520 18720
rect 24394 18708 24400 18720
rect 24452 18748 24458 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24452 18720 24593 18748
rect 24452 18708 24458 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 21508 18652 23520 18680
rect 23569 18683 23627 18689
rect 21508 18640 21514 18652
rect 23569 18649 23581 18683
rect 23615 18680 23627 18683
rect 24673 18683 24731 18689
rect 24673 18680 24685 18683
rect 23615 18652 24685 18680
rect 23615 18649 23627 18652
rect 23569 18643 23627 18649
rect 24673 18649 24685 18652
rect 24719 18649 24731 18683
rect 24780 18680 24808 18711
rect 25130 18708 25136 18760
rect 25188 18748 25194 18760
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 25188 18720 25421 18748
rect 25188 18708 25194 18720
rect 25409 18717 25421 18720
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 27338 18708 27344 18760
rect 27396 18748 27402 18760
rect 27433 18751 27491 18757
rect 27433 18748 27445 18751
rect 27396 18720 27445 18748
rect 27396 18708 27402 18720
rect 27433 18717 27445 18720
rect 27479 18717 27491 18751
rect 27433 18711 27491 18717
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28776 18720 28825 18748
rect 28776 18708 28782 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 31205 18751 31263 18757
rect 31205 18748 31217 18751
rect 28813 18711 28871 18717
rect 30300 18720 31217 18748
rect 24854 18680 24860 18692
rect 24780 18652 24860 18680
rect 24673 18643 24731 18649
rect 24854 18640 24860 18652
rect 24912 18680 24918 18692
rect 26160 18680 26188 18708
rect 30300 18692 30328 18720
rect 31205 18717 31217 18720
rect 31251 18717 31263 18751
rect 31205 18711 31263 18717
rect 31570 18708 31576 18760
rect 31628 18748 31634 18760
rect 31665 18751 31723 18757
rect 31665 18748 31677 18751
rect 31628 18720 31677 18748
rect 31628 18708 31634 18720
rect 31665 18717 31677 18720
rect 31711 18717 31723 18751
rect 31665 18711 31723 18717
rect 24912 18652 26188 18680
rect 24912 18640 24918 18652
rect 30282 18640 30288 18692
rect 30340 18640 30346 18692
rect 30926 18640 30932 18692
rect 30984 18689 30990 18692
rect 30984 18680 30996 18689
rect 30984 18652 31029 18680
rect 30984 18643 30996 18652
rect 30984 18640 30990 18643
rect 18932 18584 21041 18612
rect 18932 18572 18938 18584
rect 23382 18572 23388 18624
rect 23440 18572 23446 18624
rect 25317 18615 25375 18621
rect 25317 18581 25329 18615
rect 25363 18612 25375 18615
rect 25958 18612 25964 18624
rect 25363 18584 25964 18612
rect 25363 18581 25375 18584
rect 25317 18575 25375 18581
rect 25958 18572 25964 18584
rect 26016 18572 26022 18624
rect 29178 18572 29184 18624
rect 29236 18612 29242 18624
rect 29825 18615 29883 18621
rect 29825 18612 29837 18615
rect 29236 18584 29837 18612
rect 29236 18572 29242 18584
rect 29825 18581 29837 18584
rect 29871 18581 29883 18615
rect 29825 18575 29883 18581
rect 31757 18615 31815 18621
rect 31757 18581 31769 18615
rect 31803 18612 31815 18615
rect 32030 18612 32036 18624
rect 31803 18584 32036 18612
rect 31803 18581 31815 18584
rect 31757 18575 31815 18581
rect 32030 18572 32036 18584
rect 32088 18572 32094 18624
rect 1104 18522 32632 18544
rect 1104 18470 8792 18522
rect 8844 18470 8856 18522
rect 8908 18470 8920 18522
rect 8972 18470 8984 18522
rect 9036 18470 9048 18522
rect 9100 18470 16634 18522
rect 16686 18470 16698 18522
rect 16750 18470 16762 18522
rect 16814 18470 16826 18522
rect 16878 18470 16890 18522
rect 16942 18470 24476 18522
rect 24528 18470 24540 18522
rect 24592 18470 24604 18522
rect 24656 18470 24668 18522
rect 24720 18470 24732 18522
rect 24784 18470 32318 18522
rect 32370 18470 32382 18522
rect 32434 18470 32446 18522
rect 32498 18470 32510 18522
rect 32562 18470 32574 18522
rect 32626 18470 32632 18522
rect 1104 18448 32632 18470
rect 2590 18368 2596 18420
rect 2648 18368 2654 18420
rect 3234 18368 3240 18420
rect 3292 18408 3298 18420
rect 3697 18411 3755 18417
rect 3697 18408 3709 18411
rect 3292 18380 3709 18408
rect 3292 18368 3298 18380
rect 3697 18377 3709 18380
rect 3743 18377 3755 18411
rect 3697 18371 3755 18377
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 7167 18411 7225 18417
rect 7167 18408 7179 18411
rect 6972 18380 7179 18408
rect 6972 18368 6978 18380
rect 7167 18377 7179 18380
rect 7213 18377 7225 18411
rect 7167 18371 7225 18377
rect 8021 18411 8079 18417
rect 8021 18377 8033 18411
rect 8067 18408 8079 18411
rect 8478 18408 8484 18420
rect 8067 18380 8484 18408
rect 8067 18377 8079 18380
rect 8021 18371 8079 18377
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 9033 18411 9091 18417
rect 9033 18377 9045 18411
rect 9079 18408 9091 18411
rect 9398 18408 9404 18420
rect 9079 18380 9404 18408
rect 9079 18377 9091 18380
rect 9033 18371 9091 18377
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 10410 18368 10416 18420
rect 10468 18408 10474 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 10468 18380 10793 18408
rect 10468 18368 10474 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 12618 18368 12624 18420
rect 12676 18408 12682 18420
rect 12713 18411 12771 18417
rect 12713 18408 12725 18411
rect 12676 18380 12725 18408
rect 12676 18368 12682 18380
rect 12713 18377 12725 18380
rect 12759 18408 12771 18411
rect 12759 18380 12940 18408
rect 12759 18377 12771 18380
rect 12713 18371 12771 18377
rect 2406 18340 2412 18352
rect 2148 18312 2412 18340
rect 2148 18281 2176 18312
rect 2406 18300 2412 18312
rect 2464 18340 2470 18352
rect 5350 18340 5356 18352
rect 2464 18312 5356 18340
rect 2464 18300 2470 18312
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2363 18244 3004 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18173 2283 18207
rect 2225 18167 2283 18173
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2682 18204 2688 18216
rect 2455 18176 2688 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2240 18136 2268 18167
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 2976 18204 3004 18244
rect 3050 18232 3056 18284
rect 3108 18232 3114 18284
rect 3528 18281 3556 18312
rect 5350 18300 5356 18312
rect 5408 18300 5414 18352
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 7377 18343 7435 18349
rect 7377 18340 7389 18343
rect 7340 18312 7389 18340
rect 7340 18300 7346 18312
rect 7377 18309 7389 18312
rect 7423 18309 7435 18343
rect 8205 18343 8263 18349
rect 8205 18340 8217 18343
rect 7377 18303 7435 18309
rect 8036 18312 8217 18340
rect 8036 18284 8064 18312
rect 8205 18309 8217 18312
rect 8251 18309 8263 18343
rect 8205 18303 8263 18309
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 8849 18343 8907 18349
rect 8849 18340 8861 18343
rect 8444 18312 8861 18340
rect 8444 18300 8450 18312
rect 8849 18309 8861 18312
rect 8895 18309 8907 18343
rect 8849 18303 8907 18309
rect 8956 18312 9260 18340
rect 4430 18281 4436 18284
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 4424 18235 4436 18281
rect 4430 18232 4436 18235
rect 4488 18232 4494 18284
rect 8018 18232 8024 18284
rect 8076 18232 8082 18284
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8956 18272 8984 18312
rect 8159 18244 8984 18272
rect 9125 18275 9183 18281
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 9125 18241 9137 18275
rect 9171 18241 9183 18275
rect 9232 18272 9260 18312
rect 9950 18300 9956 18352
rect 10008 18300 10014 18352
rect 12912 18340 12940 18380
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 13688 18380 15117 18408
rect 13688 18368 13694 18380
rect 15105 18377 15117 18380
rect 15151 18377 15163 18411
rect 15105 18371 15163 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 18414 18408 18420 18420
rect 15528 18380 18420 18408
rect 15528 18368 15534 18380
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 18506 18368 18512 18420
rect 18564 18408 18570 18420
rect 19610 18408 19616 18420
rect 18564 18380 19616 18408
rect 18564 18368 18570 18380
rect 19610 18368 19616 18380
rect 19668 18408 19674 18420
rect 20254 18408 20260 18420
rect 19668 18380 20260 18408
rect 19668 18368 19674 18380
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 20346 18368 20352 18420
rect 20404 18408 20410 18420
rect 20625 18411 20683 18417
rect 20625 18408 20637 18411
rect 20404 18380 20637 18408
rect 20404 18368 20410 18380
rect 20625 18377 20637 18380
rect 20671 18377 20683 18411
rect 20625 18371 20683 18377
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 21450 18408 21456 18420
rect 21048 18380 21456 18408
rect 21048 18368 21054 18380
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 22094 18368 22100 18420
rect 22152 18368 22158 18420
rect 22738 18368 22744 18420
rect 22796 18368 22802 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 24581 18411 24639 18417
rect 24581 18408 24593 18411
rect 23440 18380 24593 18408
rect 23440 18368 23446 18380
rect 24581 18377 24593 18380
rect 24627 18377 24639 18411
rect 24581 18371 24639 18377
rect 26418 18368 26424 18420
rect 26476 18368 26482 18420
rect 18782 18340 18788 18352
rect 12912 18312 13400 18340
rect 9674 18272 9680 18284
rect 9232 18244 9680 18272
rect 9125 18235 9183 18241
rect 3326 18204 3332 18216
rect 2976 18176 3332 18204
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 4154 18164 4160 18216
rect 4212 18164 4218 18216
rect 7098 18164 7104 18216
rect 7156 18204 7162 18216
rect 7650 18204 7656 18216
rect 7156 18176 7656 18204
rect 7156 18164 7162 18176
rect 7650 18164 7656 18176
rect 7708 18204 7714 18216
rect 8128 18204 8156 18235
rect 9140 18204 9168 18235
rect 7708 18176 8156 18204
rect 8312 18176 9168 18204
rect 9646 18232 9680 18244
rect 9732 18232 9738 18284
rect 11054 18232 11060 18284
rect 11112 18232 11118 18284
rect 11146 18232 11152 18284
rect 11204 18232 11210 18284
rect 11422 18232 11428 18284
rect 11480 18272 11486 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 11480 18244 12265 18272
rect 11480 18232 11486 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12342 18232 12348 18284
rect 12400 18232 12406 18284
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 13372 18281 13400 18312
rect 13464 18312 18788 18340
rect 13464 18281 13492 18312
rect 18782 18300 18788 18312
rect 18840 18300 18846 18352
rect 20898 18340 20904 18352
rect 20088 18312 20904 18340
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 12952 18244 13185 18272
rect 12952 18232 12958 18244
rect 13173 18241 13185 18244
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18241 13415 18275
rect 13357 18235 13415 18241
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 9646 18204 9674 18232
rect 13464 18204 13492 18235
rect 14274 18232 14280 18284
rect 14332 18272 14338 18284
rect 14829 18275 14887 18281
rect 14829 18272 14841 18275
rect 14332 18244 14841 18272
rect 14332 18232 14338 18244
rect 14829 18241 14841 18244
rect 14875 18272 14887 18275
rect 14918 18272 14924 18284
rect 14875 18244 14924 18272
rect 14875 18241 14887 18244
rect 14829 18235 14887 18241
rect 14918 18232 14924 18244
rect 14976 18232 14982 18284
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18272 15163 18275
rect 15654 18272 15660 18284
rect 15151 18244 15660 18272
rect 15151 18241 15163 18244
rect 15105 18235 15163 18241
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 15470 18204 15476 18216
rect 9646 18176 13492 18204
rect 13648 18176 15476 18204
rect 7708 18164 7714 18176
rect 2148 18108 2268 18136
rect 2148 18080 2176 18108
rect 7006 18096 7012 18148
rect 7064 18096 7070 18148
rect 8312 18136 8340 18176
rect 7208 18108 8340 18136
rect 8389 18139 8447 18145
rect 7208 18080 7236 18108
rect 8389 18105 8401 18139
rect 8435 18136 8447 18139
rect 8570 18136 8576 18148
rect 8435 18108 8576 18136
rect 8435 18105 8447 18108
rect 8389 18099 8447 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8662 18096 8668 18148
rect 8720 18136 8726 18148
rect 8849 18139 8907 18145
rect 8849 18136 8861 18139
rect 8720 18108 8861 18136
rect 8720 18096 8726 18108
rect 8849 18105 8861 18108
rect 8895 18105 8907 18139
rect 12894 18136 12900 18148
rect 8849 18099 8907 18105
rect 8956 18108 12900 18136
rect 2130 18028 2136 18080
rect 2188 18028 2194 18080
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 3145 18071 3203 18077
rect 3145 18068 3157 18071
rect 2280 18040 3157 18068
rect 2280 18028 2286 18040
rect 3145 18037 3157 18040
rect 3191 18037 3203 18071
rect 3145 18031 3203 18037
rect 5537 18071 5595 18077
rect 5537 18037 5549 18071
rect 5583 18068 5595 18071
rect 6086 18068 6092 18080
rect 5583 18040 6092 18068
rect 5583 18037 5595 18040
rect 5537 18031 5595 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 7190 18028 7196 18080
rect 7248 18028 7254 18080
rect 7558 18028 7564 18080
rect 7616 18068 7622 18080
rect 7837 18071 7895 18077
rect 7837 18068 7849 18071
rect 7616 18040 7849 18068
rect 7616 18028 7622 18040
rect 7837 18037 7849 18040
rect 7883 18037 7895 18071
rect 7837 18031 7895 18037
rect 8018 18028 8024 18080
rect 8076 18068 8082 18080
rect 8956 18068 8984 18108
rect 12894 18096 12900 18108
rect 12952 18096 12958 18148
rect 13648 18145 13676 18176
rect 15470 18164 15476 18176
rect 15528 18204 15534 18216
rect 15765 18204 15793 18235
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16117 18275 16175 18281
rect 16117 18272 16129 18275
rect 15988 18244 16129 18272
rect 15988 18232 15994 18244
rect 16117 18241 16129 18244
rect 16163 18272 16175 18275
rect 20088 18272 20116 18312
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 29356 18343 29414 18349
rect 22020 18312 22692 18340
rect 22020 18284 22048 18312
rect 16163 18244 20116 18272
rect 20165 18275 20223 18281
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 20165 18241 20177 18275
rect 20211 18272 20223 18275
rect 20254 18272 20260 18284
rect 20211 18244 20260 18272
rect 20211 18241 20223 18244
rect 20165 18235 20223 18241
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 22002 18232 22008 18284
rect 22060 18232 22066 18284
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22152 18244 22201 18272
rect 22152 18232 22158 18244
rect 22189 18241 22201 18244
rect 22235 18272 22247 18275
rect 22554 18272 22560 18284
rect 22235 18244 22560 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 22664 18281 22692 18312
rect 29356 18309 29368 18343
rect 29402 18340 29414 18343
rect 31662 18340 31668 18352
rect 29402 18312 31668 18340
rect 29402 18309 29414 18312
rect 29356 18303 29414 18309
rect 31662 18300 31668 18312
rect 31720 18300 31726 18352
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18241 22707 18275
rect 22649 18235 22707 18241
rect 22738 18232 22744 18284
rect 22796 18272 22802 18284
rect 22833 18275 22891 18281
rect 22833 18272 22845 18275
rect 22796 18244 22845 18272
rect 22796 18232 22802 18244
rect 22833 18241 22845 18244
rect 22879 18241 22891 18275
rect 22833 18235 22891 18241
rect 24026 18232 24032 18284
rect 24084 18232 24090 18284
rect 24394 18232 24400 18284
rect 24452 18272 24458 18284
rect 24489 18275 24547 18281
rect 24489 18272 24501 18275
rect 24452 18244 24501 18272
rect 24452 18232 24458 18244
rect 24489 18241 24501 18244
rect 24535 18241 24547 18275
rect 24489 18235 24547 18241
rect 24673 18275 24731 18281
rect 24673 18241 24685 18275
rect 24719 18272 24731 18275
rect 24854 18272 24860 18284
rect 24719 18244 24860 18272
rect 24719 18241 24731 18244
rect 24673 18235 24731 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 26053 18275 26111 18281
rect 26053 18241 26065 18275
rect 26099 18272 26111 18275
rect 26326 18272 26332 18284
rect 26099 18244 26332 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 26326 18232 26332 18244
rect 26384 18232 26390 18284
rect 27430 18232 27436 18284
rect 27488 18232 27494 18284
rect 28077 18275 28135 18281
rect 28077 18241 28089 18275
rect 28123 18272 28135 18275
rect 29178 18272 29184 18284
rect 28123 18244 29184 18272
rect 28123 18241 28135 18244
rect 28077 18235 28135 18241
rect 29178 18232 29184 18244
rect 29236 18232 29242 18284
rect 15528 18176 15793 18204
rect 15528 18164 15534 18176
rect 19242 18164 19248 18216
rect 19300 18164 19306 18216
rect 25961 18207 26019 18213
rect 25961 18204 25973 18207
rect 19453 18176 25973 18204
rect 13633 18139 13691 18145
rect 13633 18105 13645 18139
rect 13679 18105 13691 18139
rect 13633 18099 13691 18105
rect 15010 18096 15016 18148
rect 15068 18096 15074 18148
rect 18782 18096 18788 18148
rect 18840 18136 18846 18148
rect 19453 18136 19481 18176
rect 25961 18173 25973 18176
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 29086 18164 29092 18216
rect 29144 18164 29150 18216
rect 30929 18207 30987 18213
rect 30929 18173 30941 18207
rect 30975 18173 30987 18207
rect 30929 18167 30987 18173
rect 18840 18108 19481 18136
rect 18840 18096 18846 18108
rect 19518 18096 19524 18148
rect 19576 18096 19582 18148
rect 22002 18136 22008 18148
rect 19628 18108 22008 18136
rect 8076 18040 8984 18068
rect 8076 18028 8082 18040
rect 10042 18028 10048 18080
rect 10100 18028 10106 18080
rect 11149 18071 11207 18077
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11698 18068 11704 18080
rect 11195 18040 11704 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 12492 18040 13461 18068
rect 12492 18028 12498 18040
rect 13449 18037 13461 18040
rect 13495 18068 13507 18071
rect 13722 18068 13728 18080
rect 13495 18040 13728 18068
rect 13495 18037 13507 18040
rect 13449 18031 13507 18037
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 14182 18028 14188 18080
rect 14240 18028 14246 18080
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 15286 18068 15292 18080
rect 14424 18040 15292 18068
rect 14424 18028 14430 18040
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15565 18071 15623 18077
rect 15565 18068 15577 18071
rect 15436 18040 15577 18068
rect 15436 18028 15442 18040
rect 15565 18037 15577 18040
rect 15611 18037 15623 18071
rect 15565 18031 15623 18037
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 15930 18068 15936 18080
rect 15712 18040 15936 18068
rect 15712 18028 15718 18040
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 16114 18068 16120 18080
rect 16071 18040 16120 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 16114 18028 16120 18040
rect 16172 18028 16178 18080
rect 17402 18028 17408 18080
rect 17460 18068 17466 18080
rect 19628 18068 19656 18108
rect 22002 18096 22008 18108
rect 22060 18096 22066 18148
rect 30469 18139 30527 18145
rect 30469 18105 30481 18139
rect 30515 18136 30527 18139
rect 30944 18136 30972 18167
rect 30515 18108 30972 18136
rect 30515 18105 30527 18108
rect 30469 18099 30527 18105
rect 17460 18040 19656 18068
rect 17460 18028 17466 18040
rect 19702 18028 19708 18080
rect 19760 18028 19766 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20257 18071 20315 18077
rect 20257 18068 20269 18071
rect 20220 18040 20269 18068
rect 20220 18028 20226 18040
rect 20257 18037 20269 18040
rect 20303 18037 20315 18071
rect 20257 18031 20315 18037
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 23845 18071 23903 18077
rect 23845 18068 23857 18071
rect 23440 18040 23857 18068
rect 23440 18028 23446 18040
rect 23845 18037 23857 18040
rect 23891 18037 23903 18071
rect 23845 18031 23903 18037
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 25317 18071 25375 18077
rect 25317 18068 25329 18071
rect 25280 18040 25329 18068
rect 25280 18028 25286 18040
rect 25317 18037 25329 18040
rect 25363 18037 25375 18071
rect 25317 18031 25375 18037
rect 27246 18028 27252 18080
rect 27304 18028 27310 18080
rect 28629 18071 28687 18077
rect 28629 18037 28641 18071
rect 28675 18068 28687 18071
rect 30374 18068 30380 18080
rect 28675 18040 30380 18068
rect 28675 18037 28687 18040
rect 28629 18031 28687 18037
rect 30374 18028 30380 18040
rect 30432 18028 30438 18080
rect 31570 18028 31576 18080
rect 31628 18028 31634 18080
rect 1104 17978 32476 18000
rect 1104 17926 4871 17978
rect 4923 17926 4935 17978
rect 4987 17926 4999 17978
rect 5051 17926 5063 17978
rect 5115 17926 5127 17978
rect 5179 17926 12713 17978
rect 12765 17926 12777 17978
rect 12829 17926 12841 17978
rect 12893 17926 12905 17978
rect 12957 17926 12969 17978
rect 13021 17926 20555 17978
rect 20607 17926 20619 17978
rect 20671 17926 20683 17978
rect 20735 17926 20747 17978
rect 20799 17926 20811 17978
rect 20863 17926 28397 17978
rect 28449 17926 28461 17978
rect 28513 17926 28525 17978
rect 28577 17926 28589 17978
rect 28641 17926 28653 17978
rect 28705 17926 32476 17978
rect 1104 17904 32476 17926
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2406 17864 2412 17876
rect 2363 17836 2412 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2406 17824 2412 17836
rect 2464 17824 2470 17876
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3050 17864 3056 17876
rect 3007 17836 3056 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 3602 17864 3608 17876
rect 3375 17836 3608 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 3970 17824 3976 17876
rect 4028 17864 4034 17876
rect 4028 17836 4200 17864
rect 4028 17824 4034 17836
rect 2501 17799 2559 17805
rect 2501 17765 2513 17799
rect 2547 17796 2559 17799
rect 3418 17796 3424 17808
rect 2547 17768 3424 17796
rect 2547 17765 2559 17768
rect 2501 17759 2559 17765
rect 3418 17756 3424 17768
rect 3476 17796 3482 17808
rect 4065 17799 4123 17805
rect 4065 17796 4077 17799
rect 3476 17768 4077 17796
rect 3476 17756 3482 17768
rect 4065 17765 4077 17768
rect 4111 17765 4123 17799
rect 4172 17796 4200 17836
rect 4430 17824 4436 17876
rect 4488 17824 4494 17876
rect 10042 17864 10048 17876
rect 6932 17836 10048 17864
rect 4172 17768 6408 17796
rect 4065 17759 4123 17765
rect 3142 17688 3148 17740
rect 3200 17728 3206 17740
rect 3200 17700 4200 17728
rect 3200 17688 3206 17700
rect 3050 17620 3056 17672
rect 3108 17660 3114 17672
rect 3237 17663 3295 17669
rect 3237 17660 3249 17663
rect 3108 17632 3249 17660
rect 3108 17620 3114 17632
rect 3237 17629 3249 17632
rect 3283 17629 3295 17663
rect 3237 17623 3295 17629
rect 3329 17663 3387 17669
rect 3329 17629 3341 17663
rect 3375 17629 3387 17663
rect 3329 17623 3387 17629
rect 2130 17552 2136 17604
rect 2188 17592 2194 17604
rect 2188 17564 2636 17592
rect 2188 17552 2194 17564
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2333 17527 2391 17533
rect 2333 17524 2345 17527
rect 2096 17496 2345 17524
rect 2096 17484 2102 17496
rect 2333 17493 2345 17496
rect 2379 17493 2391 17527
rect 2608 17524 2636 17564
rect 3142 17552 3148 17604
rect 3200 17592 3206 17604
rect 3344 17592 3372 17623
rect 3970 17620 3976 17672
rect 4028 17620 4034 17672
rect 4172 17669 4200 17700
rect 4172 17663 4247 17669
rect 4172 17632 4201 17663
rect 4189 17629 4201 17632
rect 4235 17629 4247 17663
rect 4189 17623 4247 17629
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 3200 17564 3372 17592
rect 3200 17552 3206 17564
rect 6086 17552 6092 17604
rect 6144 17552 6150 17604
rect 3786 17524 3792 17536
rect 2608 17496 3792 17524
rect 2333 17487 2391 17493
rect 3786 17484 3792 17496
rect 3844 17524 3850 17536
rect 5350 17524 5356 17536
rect 3844 17496 5356 17524
rect 3844 17484 3850 17496
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 6380 17533 6408 17768
rect 6932 17669 6960 17836
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 11422 17824 11428 17876
rect 11480 17824 11486 17876
rect 11974 17824 11980 17876
rect 12032 17864 12038 17876
rect 12161 17867 12219 17873
rect 12161 17864 12173 17867
rect 12032 17836 12173 17864
rect 12032 17824 12038 17836
rect 12161 17833 12173 17836
rect 12207 17833 12219 17867
rect 14734 17864 14740 17876
rect 12161 17827 12219 17833
rect 12406 17836 14740 17864
rect 7009 17799 7067 17805
rect 7009 17765 7021 17799
rect 7055 17796 7067 17799
rect 8018 17796 8024 17808
rect 7055 17768 8024 17796
rect 7055 17765 7067 17768
rect 7009 17759 7067 17765
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 10226 17796 10232 17808
rect 8352 17768 10232 17796
rect 8352 17756 8358 17768
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 10594 17756 10600 17808
rect 10652 17756 10658 17808
rect 11146 17796 11152 17808
rect 10704 17768 11152 17796
rect 10612 17728 10640 17756
rect 7116 17700 10640 17728
rect 7116 17669 7144 17700
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8386 17660 8392 17672
rect 7975 17632 8392 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8570 17620 8576 17672
rect 8628 17620 8634 17672
rect 9306 17620 9312 17672
rect 9364 17620 9370 17672
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 9858 17660 9864 17672
rect 9815 17632 9864 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 9950 17620 9956 17672
rect 10008 17620 10014 17672
rect 10597 17663 10655 17669
rect 10597 17629 10609 17663
rect 10643 17660 10655 17663
rect 10704 17660 10732 17768
rect 11146 17756 11152 17768
rect 11204 17756 11210 17808
rect 11698 17756 11704 17808
rect 11756 17756 11762 17808
rect 12406 17796 12434 17836
rect 14734 17824 14740 17836
rect 14792 17824 14798 17876
rect 15194 17864 15200 17876
rect 14927 17836 15200 17864
rect 11808 17768 12434 17796
rect 11716 17728 11744 17756
rect 10796 17700 11744 17728
rect 10796 17669 10824 17700
rect 10643 17632 10732 17660
rect 10781 17663 10839 17669
rect 10643 17629 10655 17632
rect 10597 17623 10655 17629
rect 10781 17629 10793 17663
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 11204 17632 11253 17660
rect 11204 17620 11210 17632
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 6730 17552 6736 17604
rect 6788 17592 6794 17604
rect 7558 17592 7564 17604
rect 6788 17564 7564 17592
rect 6788 17552 6794 17564
rect 7558 17552 7564 17564
rect 7616 17552 7622 17604
rect 7742 17552 7748 17604
rect 7800 17552 7806 17604
rect 8481 17595 8539 17601
rect 8481 17561 8493 17595
rect 8527 17592 8539 17595
rect 11054 17592 11060 17604
rect 8527 17564 11060 17592
rect 8527 17561 8539 17564
rect 8481 17555 8539 17561
rect 11054 17552 11060 17564
rect 11112 17552 11118 17604
rect 11256 17592 11284 17623
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 11425 17663 11483 17669
rect 11425 17660 11437 17663
rect 11388 17632 11437 17660
rect 11388 17620 11394 17632
rect 11425 17629 11437 17632
rect 11471 17629 11483 17663
rect 11425 17623 11483 17629
rect 11808 17592 11836 17768
rect 12710 17756 12716 17808
rect 12768 17796 12774 17808
rect 14366 17796 14372 17808
rect 12768 17768 14372 17796
rect 12768 17756 12774 17768
rect 14366 17756 14372 17768
rect 14424 17756 14430 17808
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 12268 17700 14749 17728
rect 12268 17650 12296 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 12345 17657 12403 17663
rect 12345 17650 12357 17657
rect 12268 17623 12357 17650
rect 12391 17623 12403 17657
rect 12268 17622 12403 17623
rect 12345 17617 12403 17622
rect 12710 17620 12716 17672
rect 12768 17620 12774 17672
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 13446 17660 13452 17672
rect 12851 17632 13452 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 11256 17564 11836 17592
rect 12434 17552 12440 17604
rect 12492 17552 12498 17604
rect 12526 17552 12532 17604
rect 12584 17552 12590 17604
rect 12820 17592 12848 17623
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17660 13599 17663
rect 14274 17660 14280 17672
rect 13587 17632 14280 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 14927 17669 14955 17836
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 19518 17864 19524 17876
rect 15344 17836 19524 17864
rect 15344 17824 15350 17836
rect 19518 17824 19524 17836
rect 19576 17864 19582 17876
rect 19886 17864 19892 17876
rect 19576 17836 19892 17864
rect 19576 17824 19582 17836
rect 19886 17824 19892 17836
rect 19944 17824 19950 17876
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 23198 17864 23204 17876
rect 20027 17836 23204 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 23477 17867 23535 17873
rect 23477 17833 23489 17867
rect 23523 17864 23535 17867
rect 23750 17864 23756 17876
rect 23523 17836 23756 17864
rect 23523 17833 23535 17836
rect 23477 17827 23535 17833
rect 23750 17824 23756 17836
rect 23808 17824 23814 17876
rect 25130 17824 25136 17876
rect 25188 17864 25194 17876
rect 31110 17864 31116 17876
rect 25188 17836 31116 17864
rect 25188 17824 25194 17836
rect 31110 17824 31116 17836
rect 31168 17824 31174 17876
rect 15013 17799 15071 17805
rect 15013 17765 15025 17799
rect 15059 17796 15071 17799
rect 19426 17796 19432 17808
rect 15059 17768 15976 17796
rect 15059 17765 15071 17768
rect 15013 17759 15071 17765
rect 15948 17728 15976 17768
rect 16132 17768 19432 17796
rect 16132 17728 16160 17768
rect 19426 17756 19432 17768
rect 19484 17756 19490 17808
rect 19702 17796 19708 17808
rect 19536 17768 19708 17796
rect 15120 17700 15516 17728
rect 15948 17700 16160 17728
rect 15120 17672 15148 17700
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15102 17620 15108 17672
rect 15160 17620 15166 17672
rect 15197 17663 15255 17669
rect 15197 17629 15209 17663
rect 15243 17662 15255 17663
rect 15243 17660 15332 17662
rect 15378 17660 15384 17672
rect 15243 17634 15384 17660
rect 15243 17629 15255 17634
rect 15304 17632 15384 17634
rect 15197 17623 15255 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15488 17660 15516 17700
rect 16206 17688 16212 17740
rect 16264 17688 16270 17740
rect 16316 17700 17356 17728
rect 16316 17672 16344 17700
rect 15933 17663 15991 17669
rect 15933 17660 15945 17663
rect 15488 17632 15945 17660
rect 15933 17629 15945 17632
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 16117 17663 16175 17669
rect 16117 17629 16129 17663
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 12636 17564 12848 17592
rect 6365 17527 6423 17533
rect 6365 17493 6377 17527
rect 6411 17524 6423 17527
rect 8294 17524 8300 17536
rect 6411 17496 8300 17524
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 9766 17484 9772 17536
rect 9824 17484 9830 17536
rect 11974 17484 11980 17536
rect 12032 17524 12038 17536
rect 12636 17524 12664 17564
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 13170 17592 13176 17604
rect 12952 17564 13176 17592
rect 12952 17552 12958 17564
rect 13170 17552 13176 17564
rect 13228 17552 13234 17604
rect 13262 17552 13268 17604
rect 13320 17592 13326 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 13320 17564 13369 17592
rect 13320 17552 13326 17564
rect 13357 17561 13369 17564
rect 13403 17561 13415 17595
rect 13357 17555 13415 17561
rect 13722 17552 13728 17604
rect 13780 17552 13786 17604
rect 15749 17595 15807 17601
rect 15749 17592 15761 17595
rect 13832 17564 15761 17592
rect 12032 17496 12664 17524
rect 12032 17484 12038 17496
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 13832 17524 13860 17564
rect 15749 17561 15761 17564
rect 15795 17561 15807 17595
rect 16132 17592 16160 17623
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 16482 17620 16488 17672
rect 16540 17620 16546 17672
rect 17328 17669 17356 17700
rect 17770 17688 17776 17740
rect 17828 17728 17834 17740
rect 19536 17737 19564 17768
rect 19702 17756 19708 17768
rect 19760 17756 19766 17808
rect 20898 17756 20904 17808
rect 20956 17796 20962 17808
rect 23566 17796 23572 17808
rect 20956 17768 23572 17796
rect 20956 17756 20962 17768
rect 23566 17756 23572 17768
rect 23624 17756 23630 17808
rect 19521 17731 19579 17737
rect 17828 17700 19288 17728
rect 17828 17688 17834 17700
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17126 17592 17132 17604
rect 16132 17564 17132 17592
rect 15749 17555 15807 17561
rect 17126 17552 17132 17564
rect 17184 17552 17190 17604
rect 17236 17592 17264 17623
rect 17402 17620 17408 17672
rect 17460 17660 17466 17672
rect 17497 17663 17555 17669
rect 17497 17660 17509 17663
rect 17460 17632 17509 17660
rect 17460 17620 17466 17632
rect 17497 17629 17509 17632
rect 17543 17629 17555 17663
rect 17497 17623 17555 17629
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 17644 17632 18368 17660
rect 17644 17620 17650 17632
rect 17236 17564 18276 17592
rect 12768 17496 13860 17524
rect 12768 17484 12774 17496
rect 17678 17484 17684 17536
rect 17736 17524 17742 17536
rect 18248 17533 18276 17564
rect 17773 17527 17831 17533
rect 17773 17524 17785 17527
rect 17736 17496 17785 17524
rect 17736 17484 17742 17496
rect 17773 17493 17785 17496
rect 17819 17493 17831 17527
rect 17773 17487 17831 17493
rect 18233 17527 18291 17533
rect 18233 17493 18245 17527
rect 18279 17493 18291 17527
rect 18340 17524 18368 17632
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 18472 17632 18514 17660
rect 18472 17620 18478 17632
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 18874 17620 18880 17672
rect 18932 17620 18938 17672
rect 19260 17660 19288 17700
rect 19521 17697 19533 17731
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 21082 17728 21088 17740
rect 19659 17700 21088 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 19628 17660 19656 17691
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 23106 17688 23112 17740
rect 23164 17728 23170 17740
rect 26510 17728 26516 17740
rect 23164 17700 26516 17728
rect 23164 17688 23170 17700
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 19260 17632 19656 17660
rect 19702 17620 19708 17672
rect 19760 17620 19766 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17660 19855 17663
rect 20254 17660 20260 17672
rect 19843 17632 20260 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23385 17663 23443 17669
rect 23385 17629 23397 17663
rect 23431 17660 23443 17663
rect 24854 17660 24860 17672
rect 23431 17632 24860 17660
rect 23431 17629 23443 17632
rect 23385 17623 23443 17629
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 26050 17620 26056 17672
rect 26108 17660 26114 17672
rect 28629 17663 28687 17669
rect 26108 17632 26924 17660
rect 26108 17620 26114 17632
rect 19242 17552 19248 17604
rect 19300 17592 19306 17604
rect 20714 17592 20720 17604
rect 19300 17564 20720 17592
rect 19300 17552 19306 17564
rect 20714 17552 20720 17564
rect 20772 17552 20778 17604
rect 21082 17552 21088 17604
rect 21140 17592 21146 17604
rect 23474 17592 23480 17604
rect 21140 17564 23480 17592
rect 21140 17552 21146 17564
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 23569 17595 23627 17601
rect 23569 17561 23581 17595
rect 23615 17592 23627 17595
rect 23658 17592 23664 17604
rect 23615 17564 23664 17592
rect 23615 17561 23627 17564
rect 23569 17555 23627 17561
rect 23658 17552 23664 17564
rect 23716 17592 23722 17604
rect 23716 17564 24900 17592
rect 23716 17552 23722 17564
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 18340 17496 18429 17524
rect 18233 17487 18291 17493
rect 18417 17493 18429 17496
rect 18463 17524 18475 17527
rect 19334 17524 19340 17536
rect 18463 17496 19340 17524
rect 18463 17493 18475 17496
rect 18417 17487 18475 17493
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 23109 17527 23167 17533
rect 23109 17524 23121 17527
rect 20036 17496 23121 17524
rect 20036 17484 20042 17496
rect 23109 17493 23121 17496
rect 23155 17493 23167 17527
rect 23109 17487 23167 17493
rect 23290 17484 23296 17536
rect 23348 17524 23354 17536
rect 24302 17524 24308 17536
rect 23348 17496 24308 17524
rect 23348 17484 23354 17496
rect 24302 17484 24308 17496
rect 24360 17524 24366 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24360 17496 24685 17524
rect 24360 17484 24366 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24872 17524 24900 17564
rect 24946 17552 24952 17604
rect 25004 17552 25010 17604
rect 26602 17552 26608 17604
rect 26660 17592 26666 17604
rect 26758 17595 26816 17601
rect 26758 17592 26770 17595
rect 26660 17564 26770 17592
rect 26660 17552 26666 17564
rect 26758 17561 26770 17564
rect 26804 17561 26816 17595
rect 26896 17592 26924 17632
rect 28629 17629 28641 17663
rect 28675 17660 28687 17663
rect 28718 17660 28724 17672
rect 28675 17632 28724 17660
rect 28675 17629 28687 17632
rect 28629 17623 28687 17629
rect 28718 17620 28724 17632
rect 28776 17620 28782 17672
rect 30282 17620 30288 17672
rect 30340 17660 30346 17672
rect 31297 17663 31355 17669
rect 31297 17660 31309 17663
rect 30340 17632 31309 17660
rect 30340 17620 30346 17632
rect 31297 17629 31309 17632
rect 31343 17629 31355 17663
rect 31297 17623 31355 17629
rect 31757 17663 31815 17669
rect 31757 17629 31769 17663
rect 31803 17660 31815 17663
rect 31846 17660 31852 17672
rect 31803 17632 31852 17660
rect 31803 17629 31815 17632
rect 31757 17623 31815 17629
rect 31846 17620 31852 17632
rect 31904 17620 31910 17672
rect 29730 17592 29736 17604
rect 26896 17564 29736 17592
rect 26758 17555 26816 17561
rect 29730 17552 29736 17564
rect 29788 17552 29794 17604
rect 31052 17595 31110 17601
rect 31052 17561 31064 17595
rect 31098 17592 31110 17595
rect 31570 17592 31576 17604
rect 31098 17564 31576 17592
rect 31098 17561 31110 17564
rect 31052 17555 31110 17561
rect 31570 17552 31576 17564
rect 31628 17552 31634 17604
rect 25774 17524 25780 17536
rect 24872 17496 25780 17524
rect 24673 17487 24731 17493
rect 25774 17484 25780 17496
rect 25832 17524 25838 17536
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25832 17496 25881 17524
rect 25832 17484 25838 17496
rect 25869 17493 25881 17496
rect 25915 17493 25927 17527
rect 25869 17487 25927 17493
rect 26234 17484 26240 17536
rect 26292 17524 26298 17536
rect 27430 17524 27436 17536
rect 26292 17496 27436 17524
rect 26292 17484 26298 17496
rect 27430 17484 27436 17496
rect 27488 17524 27494 17536
rect 27893 17527 27951 17533
rect 27893 17524 27905 17527
rect 27488 17496 27905 17524
rect 27488 17484 27494 17496
rect 27893 17493 27905 17496
rect 27939 17493 27951 17527
rect 27893 17487 27951 17493
rect 28813 17527 28871 17533
rect 28813 17493 28825 17527
rect 28859 17524 28871 17527
rect 29822 17524 29828 17536
rect 28859 17496 29828 17524
rect 28859 17493 28871 17496
rect 28813 17487 28871 17493
rect 29822 17484 29828 17496
rect 29880 17484 29886 17536
rect 29914 17484 29920 17536
rect 29972 17484 29978 17536
rect 30006 17484 30012 17536
rect 30064 17524 30070 17536
rect 31846 17524 31852 17536
rect 30064 17496 31852 17524
rect 30064 17484 30070 17496
rect 31846 17484 31852 17496
rect 31904 17524 31910 17536
rect 31941 17527 31999 17533
rect 31941 17524 31953 17527
rect 31904 17496 31953 17524
rect 31904 17484 31910 17496
rect 31941 17493 31953 17496
rect 31987 17493 31999 17527
rect 31941 17487 31999 17493
rect 1104 17434 32632 17456
rect 1104 17382 8792 17434
rect 8844 17382 8856 17434
rect 8908 17382 8920 17434
rect 8972 17382 8984 17434
rect 9036 17382 9048 17434
rect 9100 17382 16634 17434
rect 16686 17382 16698 17434
rect 16750 17382 16762 17434
rect 16814 17382 16826 17434
rect 16878 17382 16890 17434
rect 16942 17382 24476 17434
rect 24528 17382 24540 17434
rect 24592 17382 24604 17434
rect 24656 17382 24668 17434
rect 24720 17382 24732 17434
rect 24784 17382 32318 17434
rect 32370 17382 32382 17434
rect 32434 17382 32446 17434
rect 32498 17382 32510 17434
rect 32562 17382 32574 17434
rect 32626 17382 32632 17434
rect 1104 17360 32632 17382
rect 3326 17280 3332 17332
rect 3384 17280 3390 17332
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 3602 17320 3608 17332
rect 3476 17292 3608 17320
rect 3476 17280 3482 17292
rect 3602 17280 3608 17292
rect 3660 17320 3666 17332
rect 5445 17323 5503 17329
rect 3660 17292 4660 17320
rect 3660 17280 3666 17292
rect 2961 17255 3019 17261
rect 2961 17221 2973 17255
rect 3007 17252 3019 17255
rect 3050 17252 3056 17264
rect 3007 17224 3056 17252
rect 3007 17221 3019 17224
rect 2961 17215 3019 17221
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 3191 17221 3249 17227
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2682 17184 2688 17196
rect 2363 17156 2688 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2682 17144 2688 17156
rect 2740 17184 2746 17196
rect 3191 17187 3203 17221
rect 3237 17196 3249 17221
rect 3237 17187 3240 17196
rect 2740 17144 2774 17184
rect 3191 17181 3240 17187
rect 3192 17156 3240 17181
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4154 17184 4160 17196
rect 4111 17156 4160 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4338 17193 4344 17196
rect 4332 17147 4344 17193
rect 4338 17144 4344 17147
rect 4396 17144 4402 17196
rect 4632 17184 4660 17292
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5534 17320 5540 17332
rect 5491 17292 5540 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5460 17252 5488 17283
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 8202 17320 8208 17332
rect 6963 17292 8208 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 9493 17323 9551 17329
rect 8312 17292 9260 17320
rect 6825 17255 6883 17261
rect 6825 17252 6837 17255
rect 5460 17224 6837 17252
rect 6825 17221 6837 17224
rect 6871 17221 6883 17255
rect 6825 17215 6883 17221
rect 7006 17212 7012 17264
rect 7064 17252 7070 17264
rect 8312 17252 8340 17292
rect 7064 17224 8340 17252
rect 8380 17255 8438 17261
rect 7064 17212 7070 17224
rect 8380 17221 8392 17255
rect 8426 17252 8438 17255
rect 9122 17252 9128 17264
rect 8426 17224 9128 17252
rect 8426 17221 8438 17224
rect 8380 17215 8438 17221
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 9232 17252 9260 17292
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 9858 17320 9864 17332
rect 9539 17292 9864 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 9858 17280 9864 17292
rect 9916 17320 9922 17332
rect 12526 17320 12532 17332
rect 9916 17292 10548 17320
rect 9916 17280 9922 17292
rect 9674 17252 9680 17264
rect 9232 17224 9680 17252
rect 9674 17212 9680 17224
rect 9732 17212 9738 17264
rect 9950 17212 9956 17264
rect 10008 17252 10014 17264
rect 10134 17252 10140 17264
rect 10008 17224 10140 17252
rect 10008 17212 10014 17224
rect 10134 17212 10140 17224
rect 10192 17252 10198 17264
rect 10413 17255 10471 17261
rect 10413 17252 10425 17255
rect 10192 17224 10425 17252
rect 10192 17212 10198 17224
rect 10413 17221 10425 17224
rect 10459 17221 10471 17255
rect 10413 17215 10471 17221
rect 5994 17184 6000 17196
rect 4632 17156 6000 17184
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6086 17144 6092 17196
rect 6144 17184 6150 17196
rect 9858 17184 9864 17196
rect 6144 17182 6868 17184
rect 7015 17182 9864 17184
rect 6144 17156 9864 17182
rect 6144 17144 6150 17156
rect 6840 17154 7043 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 10520 17184 10548 17292
rect 12360 17292 12532 17320
rect 11238 17252 11244 17264
rect 10796 17224 11244 17252
rect 10796 17184 10824 17224
rect 11238 17212 11244 17224
rect 11296 17252 11302 17264
rect 11790 17252 11796 17264
rect 11296 17224 11796 17252
rect 11296 17212 11302 17224
rect 11790 17212 11796 17224
rect 11848 17212 11854 17264
rect 12360 17261 12388 17292
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 12710 17280 12716 17332
rect 12768 17280 12774 17332
rect 12894 17280 12900 17332
rect 12952 17280 12958 17332
rect 13909 17323 13967 17329
rect 13909 17320 13921 17323
rect 13195 17292 13921 17320
rect 12345 17255 12403 17261
rect 12345 17221 12357 17255
rect 12391 17221 12403 17255
rect 12345 17215 12403 17221
rect 12621 17255 12679 17261
rect 12621 17221 12633 17255
rect 12667 17252 12679 17255
rect 13195 17252 13223 17292
rect 13909 17289 13921 17292
rect 13955 17289 13967 17323
rect 13909 17283 13967 17289
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 16482 17320 16488 17332
rect 15795 17292 16488 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 17126 17280 17132 17332
rect 17184 17320 17190 17332
rect 18325 17323 18383 17329
rect 18325 17320 18337 17323
rect 17184 17292 18337 17320
rect 17184 17280 17190 17292
rect 18325 17289 18337 17292
rect 18371 17289 18383 17323
rect 18325 17283 18383 17289
rect 18693 17323 18751 17329
rect 18693 17289 18705 17323
rect 18739 17320 18751 17323
rect 19518 17320 19524 17332
rect 18739 17292 19524 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 19518 17280 19524 17292
rect 19576 17280 19582 17332
rect 19794 17280 19800 17332
rect 19852 17280 19858 17332
rect 20254 17280 20260 17332
rect 20312 17280 20318 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 23532 17292 25053 17320
rect 23532 17280 23538 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25041 17283 25099 17289
rect 26050 17280 26056 17332
rect 26108 17280 26114 17332
rect 26234 17320 26240 17332
rect 26160 17292 26240 17320
rect 17770 17252 17776 17264
rect 12667 17224 13223 17252
rect 16040 17224 17776 17252
rect 12667 17221 12679 17224
rect 12621 17215 12679 17221
rect 10275 17156 10824 17184
rect 10873 17187 10931 17193
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17085 2559 17119
rect 2746 17116 2774 17144
rect 2746 17088 4108 17116
rect 2501 17079 2559 17085
rect 2516 17048 2544 17079
rect 3326 17048 3332 17060
rect 2516 17020 3332 17048
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 2133 16983 2191 16989
rect 2133 16980 2145 16983
rect 2096 16952 2145 16980
rect 2096 16940 2102 16952
rect 2133 16949 2145 16952
rect 2179 16949 2191 16983
rect 2133 16943 2191 16949
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 3145 16983 3203 16989
rect 3145 16980 3157 16983
rect 3108 16952 3157 16980
rect 3108 16940 3114 16952
rect 3145 16949 3157 16952
rect 3191 16980 3203 16983
rect 3418 16980 3424 16992
rect 3191 16952 3424 16980
rect 3191 16949 3203 16952
rect 3145 16943 3203 16949
rect 3418 16940 3424 16952
rect 3476 16940 3482 16992
rect 4080 16980 4108 17088
rect 7098 17076 7104 17128
rect 7156 17076 7162 17128
rect 7190 17076 7196 17128
rect 7248 17076 7254 17128
rect 8110 17076 8116 17128
rect 8168 17076 8174 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 10888 17116 10916 17147
rect 11054 17144 11060 17196
rect 11112 17144 11118 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17184 11759 17187
rect 12250 17184 12256 17196
rect 11747 17156 12256 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 9824 17088 10916 17116
rect 9824 17076 9830 17088
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 5408 17020 7236 17048
rect 5408 17008 5414 17020
rect 6730 16980 6736 16992
rect 4080 16952 6736 16980
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 7006 16940 7012 16992
rect 7064 16940 7070 16992
rect 7208 16980 7236 17020
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 11716 17048 11744 17147
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 12526 17144 12532 17196
rect 12584 17144 12590 17196
rect 13354 17144 13360 17196
rect 13412 17144 13418 17196
rect 13446 17144 13452 17196
rect 13504 17144 13510 17196
rect 13630 17144 13636 17196
rect 13688 17144 13694 17196
rect 13733 17187 13791 17193
rect 13733 17153 13745 17187
rect 13779 17153 13791 17187
rect 13733 17147 13791 17153
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17116 11851 17119
rect 13740 17116 13768 17147
rect 14734 17144 14740 17196
rect 14792 17144 14798 17196
rect 16040 17193 16068 17224
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 19978 17252 19984 17264
rect 17880 17224 19984 17252
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 14844 17156 15945 17184
rect 11839 17088 13768 17116
rect 11839 17085 11851 17088
rect 11793 17079 11851 17085
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 14844 17116 14872 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 14516 17088 14872 17116
rect 15013 17119 15071 17125
rect 14516 17076 14522 17088
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 16114 17116 16120 17128
rect 15013 17079 15071 17085
rect 15304 17088 16120 17116
rect 9732 17020 11744 17048
rect 9732 17008 9738 17020
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 13630 17048 13636 17060
rect 12216 17020 13636 17048
rect 12216 17008 12222 17020
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 13722 17008 13728 17060
rect 13780 17048 13786 17060
rect 15028 17048 15056 17079
rect 15304 17057 15332 17088
rect 16114 17076 16120 17088
rect 16172 17116 16178 17128
rect 16224 17116 16252 17147
rect 16172 17088 16252 17116
rect 16172 17076 16178 17088
rect 13780 17020 15056 17048
rect 15289 17051 15347 17057
rect 13780 17008 13786 17020
rect 15289 17017 15301 17051
rect 15335 17017 15347 17051
rect 16316 17048 16344 17147
rect 17678 17144 17684 17196
rect 17736 17144 17742 17196
rect 17880 17193 17908 17224
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 23382 17261 23388 17264
rect 23376 17252 23388 17261
rect 23343 17224 23388 17252
rect 23376 17215 23388 17224
rect 23382 17212 23388 17215
rect 23440 17212 23446 17264
rect 26068 17252 26096 17280
rect 23492 17224 26096 17252
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 18506 17144 18512 17196
rect 18564 17144 18570 17196
rect 18785 17187 18843 17193
rect 18785 17153 18797 17187
rect 18831 17153 18843 17187
rect 18785 17147 18843 17153
rect 18800 17048 18828 17147
rect 19426 17144 19432 17196
rect 19484 17144 19490 17196
rect 20714 17144 20720 17196
rect 20772 17144 20778 17196
rect 21266 17144 21272 17196
rect 21324 17144 21330 17196
rect 21358 17144 21364 17196
rect 21416 17184 21422 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21416 17156 22017 17184
rect 21416 17144 21422 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22186 17144 22192 17196
rect 22244 17144 22250 17196
rect 23492 17184 23520 17224
rect 23032 17156 23520 17184
rect 19334 17076 19340 17128
rect 19392 17076 19398 17128
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 23032 17116 23060 17156
rect 24762 17144 24768 17196
rect 24820 17184 24826 17196
rect 25225 17187 25283 17193
rect 25225 17184 25237 17187
rect 24820 17156 25237 17184
rect 24820 17144 24826 17156
rect 25225 17153 25237 17156
rect 25271 17153 25283 17187
rect 25225 17147 25283 17153
rect 25498 17144 25504 17196
rect 25556 17144 25562 17196
rect 25590 17144 25596 17196
rect 25648 17184 25654 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 25648 17156 26065 17184
rect 25648 17144 25654 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 19576 17088 21404 17116
rect 19576 17076 19582 17088
rect 19978 17048 19984 17060
rect 16316 17020 18736 17048
rect 18800 17020 19984 17048
rect 15289 17011 15347 17017
rect 9398 16980 9404 16992
rect 7208 16952 9404 16980
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10042 16940 10048 16992
rect 10100 16940 10106 16992
rect 10962 16940 10968 16992
rect 11020 16940 11026 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 12618 16980 12624 16992
rect 11848 16952 12624 16980
rect 11848 16940 11854 16952
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 15068 16952 15117 16980
rect 15068 16940 15074 16952
rect 15105 16949 15117 16952
rect 15151 16980 15163 16983
rect 16022 16980 16028 16992
rect 15151 16952 16028 16980
rect 15151 16949 15163 16952
rect 15105 16943 15163 16949
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 17770 16940 17776 16992
rect 17828 16940 17834 16992
rect 18708 16980 18736 17020
rect 19978 17008 19984 17020
rect 20036 17008 20042 17060
rect 21376 17057 21404 17088
rect 21560 17088 23060 17116
rect 21361 17051 21419 17057
rect 21361 17017 21373 17051
rect 21407 17048 21419 17051
rect 21450 17048 21456 17060
rect 21407 17020 21456 17048
rect 21407 17017 21419 17020
rect 21361 17011 21419 17017
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 19794 16980 19800 16992
rect 18708 16952 19800 16980
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 19944 16952 20453 16980
rect 19944 16940 19950 16952
rect 20441 16949 20453 16952
rect 20487 16949 20499 16983
rect 20441 16943 20499 16949
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 21560 16980 21588 17088
rect 23106 17076 23112 17128
rect 23164 17076 23170 17128
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17116 25467 17119
rect 26160 17116 26188 17292
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 26326 17280 26332 17332
rect 26384 17280 26390 17332
rect 26602 17280 26608 17332
rect 26660 17280 26666 17332
rect 26344 17252 26372 17280
rect 29549 17255 29607 17261
rect 29549 17252 29561 17255
rect 26344 17224 29561 17252
rect 29549 17221 29561 17224
rect 29595 17221 29607 17255
rect 29549 17215 29607 17221
rect 30374 17212 30380 17264
rect 30432 17252 30438 17264
rect 30530 17255 30588 17261
rect 30530 17252 30542 17255
rect 30432 17224 30542 17252
rect 30432 17212 30438 17224
rect 30530 17221 30542 17224
rect 30576 17221 30588 17255
rect 30530 17215 30588 17221
rect 26234 17144 26240 17196
rect 26292 17144 26298 17196
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 26344 17116 26372 17147
rect 26418 17144 26424 17196
rect 26476 17144 26482 17196
rect 28258 17144 28264 17196
rect 28316 17184 28322 17196
rect 28546 17187 28604 17193
rect 28546 17184 28558 17187
rect 28316 17156 28558 17184
rect 28316 17144 28322 17156
rect 28546 17153 28558 17156
rect 28592 17153 28604 17187
rect 28546 17147 28604 17153
rect 29825 17187 29883 17193
rect 29825 17153 29837 17187
rect 29871 17184 29883 17187
rect 30006 17184 30012 17196
rect 29871 17156 30012 17184
rect 29871 17153 29883 17156
rect 29825 17147 29883 17153
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 27246 17116 27252 17128
rect 25455 17088 26188 17116
rect 26252 17088 27252 17116
rect 25455 17085 25467 17088
rect 25409 17079 25467 17085
rect 24489 17051 24547 17057
rect 24489 17017 24501 17051
rect 24535 17048 24547 17051
rect 24946 17048 24952 17060
rect 24535 17020 24952 17048
rect 24535 17017 24547 17020
rect 24489 17011 24547 17017
rect 24946 17008 24952 17020
rect 25004 17048 25010 17060
rect 25004 17020 25268 17048
rect 25004 17008 25010 17020
rect 20772 16952 21588 16980
rect 22005 16983 22063 16989
rect 20772 16940 20778 16952
rect 22005 16949 22017 16983
rect 22051 16980 22063 16983
rect 22094 16980 22100 16992
rect 22051 16952 22100 16980
rect 22051 16949 22063 16952
rect 22005 16943 22063 16949
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 25240 16989 25268 17020
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 26252 17048 26280 17088
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 28810 17076 28816 17128
rect 28868 17076 28874 17128
rect 29086 17076 29092 17128
rect 29144 17116 29150 17128
rect 30282 17116 30288 17128
rect 29144 17088 30288 17116
rect 29144 17076 29150 17088
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 25740 17020 26280 17048
rect 27264 17048 27292 17076
rect 27264 17020 27936 17048
rect 25740 17008 25746 17020
rect 25225 16983 25283 16989
rect 25225 16949 25237 16983
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 25498 16940 25504 16992
rect 25556 16980 25562 16992
rect 26142 16980 26148 16992
rect 25556 16952 26148 16980
rect 25556 16940 25562 16952
rect 26142 16940 26148 16952
rect 26200 16980 26206 16992
rect 27433 16983 27491 16989
rect 27433 16980 27445 16983
rect 26200 16952 27445 16980
rect 26200 16940 26206 16952
rect 27433 16949 27445 16952
rect 27479 16980 27491 16983
rect 27614 16980 27620 16992
rect 27479 16952 27620 16980
rect 27479 16949 27491 16952
rect 27433 16943 27491 16949
rect 27614 16940 27620 16952
rect 27672 16940 27678 16992
rect 27908 16980 27936 17020
rect 28902 16980 28908 16992
rect 27908 16952 28908 16980
rect 28902 16940 28908 16952
rect 28960 16940 28966 16992
rect 30466 16940 30472 16992
rect 30524 16980 30530 16992
rect 31665 16983 31723 16989
rect 31665 16980 31677 16983
rect 30524 16952 31677 16980
rect 30524 16940 30530 16952
rect 31665 16949 31677 16952
rect 31711 16949 31723 16983
rect 31665 16943 31723 16949
rect 1104 16890 32476 16912
rect 1104 16838 4871 16890
rect 4923 16838 4935 16890
rect 4987 16838 4999 16890
rect 5051 16838 5063 16890
rect 5115 16838 5127 16890
rect 5179 16838 12713 16890
rect 12765 16838 12777 16890
rect 12829 16838 12841 16890
rect 12893 16838 12905 16890
rect 12957 16838 12969 16890
rect 13021 16838 20555 16890
rect 20607 16838 20619 16890
rect 20671 16838 20683 16890
rect 20735 16838 20747 16890
rect 20799 16838 20811 16890
rect 20863 16838 28397 16890
rect 28449 16838 28461 16890
rect 28513 16838 28525 16890
rect 28577 16838 28589 16890
rect 28641 16838 28653 16890
rect 28705 16838 32476 16890
rect 1104 16816 32476 16838
rect 4154 16776 4160 16788
rect 3988 16748 4160 16776
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 2038 16532 2044 16584
rect 2096 16532 2102 16584
rect 2130 16532 2136 16584
rect 2188 16532 2194 16584
rect 2332 16572 2360 16671
rect 2682 16600 2688 16652
rect 2740 16640 2746 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2740 16612 2973 16640
rect 2740 16600 2746 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3050 16600 3056 16652
rect 3108 16600 3114 16652
rect 3142 16600 3148 16652
rect 3200 16600 3206 16652
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3988 16649 4016 16748
rect 4154 16736 4160 16748
rect 4212 16776 4218 16788
rect 8110 16776 8116 16788
rect 4212 16748 8116 16776
rect 4212 16736 4218 16748
rect 5920 16649 5948 16748
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16776 8447 16779
rect 10042 16776 10048 16788
rect 8435 16748 10048 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 12529 16779 12587 16785
rect 12529 16776 12541 16779
rect 12492 16748 12541 16776
rect 12492 16736 12498 16748
rect 12529 16745 12541 16748
rect 12575 16745 12587 16779
rect 12529 16739 12587 16745
rect 14550 16736 14556 16788
rect 14608 16736 14614 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14792 16748 15025 16776
rect 14792 16736 14798 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 15933 16779 15991 16785
rect 15933 16776 15945 16779
rect 15804 16748 15945 16776
rect 15804 16736 15810 16748
rect 15933 16745 15945 16748
rect 15979 16745 15991 16779
rect 15933 16739 15991 16745
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16080 16748 20300 16776
rect 16080 16736 16086 16748
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 7248 16680 7297 16708
rect 7248 16668 7254 16680
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 7285 16671 7343 16677
rect 8573 16711 8631 16717
rect 8573 16677 8585 16711
rect 8619 16708 8631 16711
rect 9306 16708 9312 16720
rect 8619 16680 9312 16708
rect 8619 16677 8631 16680
rect 8573 16671 8631 16677
rect 3973 16643 4031 16649
rect 3292 16612 3924 16640
rect 3292 16600 3298 16612
rect 3160 16572 3188 16600
rect 3602 16572 3608 16584
rect 2332 16544 3004 16572
rect 3160 16544 3608 16572
rect 2314 16464 2320 16516
rect 2372 16464 2378 16516
rect 2777 16439 2835 16445
rect 2777 16405 2789 16439
rect 2823 16436 2835 16439
rect 2866 16436 2872 16448
rect 2823 16408 2872 16436
rect 2823 16405 2835 16408
rect 2777 16399 2835 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 2976 16436 3004 16544
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 3896 16572 3924 16612
rect 3973 16609 3985 16643
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16609 5963 16643
rect 7300 16640 7328 16671
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 9398 16668 9404 16720
rect 9456 16708 9462 16720
rect 12618 16708 12624 16720
rect 9456 16680 12624 16708
rect 9456 16668 9462 16680
rect 8202 16640 8208 16652
rect 7300 16612 8208 16640
rect 5905 16603 5963 16609
rect 8202 16600 8208 16612
rect 8260 16640 8266 16652
rect 9585 16643 9643 16649
rect 9585 16640 9597 16643
rect 8260 16612 9597 16640
rect 8260 16600 8266 16612
rect 9585 16609 9597 16612
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9674 16600 9680 16652
rect 9732 16600 9738 16652
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 10226 16640 10232 16652
rect 9815 16612 10232 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10410 16600 10416 16652
rect 10468 16600 10474 16652
rect 10888 16649 10916 16680
rect 12618 16668 12624 16680
rect 12676 16708 12682 16720
rect 12805 16711 12863 16717
rect 12805 16708 12817 16711
rect 12676 16680 12817 16708
rect 12676 16668 12682 16680
rect 12805 16677 12817 16680
rect 12851 16708 12863 16711
rect 13446 16708 13452 16720
rect 12851 16680 13452 16708
rect 12851 16677 12863 16680
rect 12805 16671 12863 16677
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 14826 16668 14832 16720
rect 14884 16708 14890 16720
rect 16393 16711 16451 16717
rect 16393 16708 16405 16711
rect 14884 16680 16405 16708
rect 14884 16668 14890 16680
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16609 10931 16643
rect 10873 16603 10931 16609
rect 11422 16600 11428 16652
rect 11480 16640 11486 16652
rect 12897 16643 12955 16649
rect 11480 16612 12112 16640
rect 11480 16600 11486 16612
rect 9493 16575 9551 16581
rect 3896 16544 4936 16572
rect 4246 16513 4252 16516
rect 4240 16467 4252 16513
rect 4246 16464 4252 16467
rect 4304 16464 4310 16516
rect 4338 16436 4344 16448
rect 2976 16408 4344 16436
rect 4338 16396 4344 16408
rect 4396 16396 4402 16448
rect 4908 16436 4936 16544
rect 9493 16541 9505 16575
rect 9539 16572 9551 16575
rect 9539 16544 9674 16572
rect 9539 16541 9551 16544
rect 9493 16535 9551 16541
rect 5258 16464 5264 16516
rect 5316 16504 5322 16516
rect 6150 16507 6208 16513
rect 6150 16504 6162 16507
rect 5316 16476 6162 16504
rect 5316 16464 5322 16476
rect 6150 16473 6162 16476
rect 6196 16473 6208 16507
rect 6150 16467 6208 16473
rect 7282 16464 7288 16516
rect 7340 16504 7346 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 7340 16476 8217 16504
rect 7340 16464 7346 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 9646 16504 9674 16544
rect 9950 16532 9956 16584
rect 10008 16572 10014 16584
rect 10597 16575 10655 16581
rect 10597 16572 10609 16575
rect 10008 16544 10609 16572
rect 10008 16532 10014 16544
rect 10597 16541 10609 16544
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 10410 16504 10416 16516
rect 9646 16476 10416 16504
rect 8205 16467 8263 16473
rect 10410 16464 10416 16476
rect 10468 16464 10474 16516
rect 10612 16504 10640 16535
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 11606 16572 11612 16584
rect 10836 16544 11612 16572
rect 10836 16532 10842 16544
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 11882 16532 11888 16584
rect 11940 16532 11946 16584
rect 12084 16581 12112 16612
rect 12897 16609 12909 16643
rect 12943 16640 12955 16643
rect 13354 16640 13360 16652
rect 12943 16612 13360 16640
rect 12943 16609 12955 16612
rect 12897 16603 12955 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 14424 16612 14657 16640
rect 14424 16600 14430 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15160 16612 15485 16640
rect 15160 16600 15166 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15672 16640 15700 16680
rect 16393 16677 16405 16680
rect 16439 16677 16451 16711
rect 20272 16708 20300 16748
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 21361 16779 21419 16785
rect 21361 16776 21373 16779
rect 20956 16748 21373 16776
rect 20956 16736 20962 16748
rect 21361 16745 21373 16748
rect 21407 16745 21419 16779
rect 23106 16776 23112 16788
rect 21361 16739 21419 16745
rect 22020 16748 23112 16776
rect 21082 16708 21088 16720
rect 20272 16680 21088 16708
rect 16393 16671 16451 16677
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 15672 16612 15792 16640
rect 15473 16603 15531 16609
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12713 16575 12771 16581
rect 12713 16572 12725 16575
rect 12308 16544 12725 16572
rect 12308 16532 12314 16544
rect 12713 16541 12725 16544
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 12986 16532 12992 16584
rect 13044 16532 13050 16584
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16572 13231 16575
rect 13446 16572 13452 16584
rect 13219 16544 13452 16572
rect 13219 16541 13231 16544
rect 13173 16535 13231 16541
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 14826 16532 14832 16584
rect 14884 16532 14890 16584
rect 15565 16575 15623 16581
rect 15565 16541 15577 16575
rect 15611 16572 15623 16575
rect 15654 16572 15660 16584
rect 15611 16544 15660 16572
rect 15611 16541 15623 16544
rect 15565 16535 15623 16541
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 15764 16581 15792 16612
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 19484 16612 20177 16640
rect 19484 16600 19490 16612
rect 20165 16609 20177 16612
rect 20211 16640 20223 16643
rect 21266 16640 21272 16652
rect 20211 16612 21272 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 21266 16600 21272 16612
rect 21324 16640 21330 16652
rect 21910 16640 21916 16652
rect 21324 16612 21916 16640
rect 21324 16600 21330 16612
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 22020 16649 22048 16748
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 24360 16748 24777 16776
rect 24360 16736 24366 16748
rect 24765 16745 24777 16748
rect 24811 16745 24823 16779
rect 25222 16776 25228 16788
rect 24765 16739 24823 16745
rect 24872 16748 25228 16776
rect 24872 16708 24900 16748
rect 25222 16736 25228 16748
rect 25280 16736 25286 16788
rect 26510 16736 26516 16788
rect 26568 16776 26574 16788
rect 27341 16779 27399 16785
rect 27341 16776 27353 16779
rect 26568 16748 27353 16776
rect 26568 16736 26574 16748
rect 27341 16745 27353 16748
rect 27387 16776 27399 16779
rect 29086 16776 29092 16788
rect 27387 16748 29092 16776
rect 27387 16745 27399 16748
rect 27341 16739 27399 16745
rect 29086 16736 29092 16748
rect 29144 16736 29150 16788
rect 31110 16736 31116 16788
rect 31168 16736 31174 16788
rect 23768 16680 24900 16708
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 16390 16532 16396 16584
rect 16448 16532 16454 16584
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 17497 16575 17555 16581
rect 17497 16572 17509 16575
rect 16540 16544 17509 16572
rect 16540 16532 16546 16544
rect 17497 16541 17509 16544
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 19702 16572 19708 16584
rect 17727 16544 19708 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19978 16532 19984 16584
rect 20036 16532 20042 16584
rect 21008 16544 22048 16572
rect 21008 16516 21036 16544
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 10612 16476 14565 16504
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 16669 16507 16727 16513
rect 16669 16504 16681 16507
rect 15988 16476 16681 16504
rect 15988 16464 15994 16476
rect 16669 16473 16681 16476
rect 16715 16504 16727 16507
rect 19426 16504 19432 16516
rect 16715 16476 19432 16504
rect 16715 16473 16727 16476
rect 16669 16467 16727 16473
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 19794 16464 19800 16516
rect 19852 16504 19858 16516
rect 19852 16476 20024 16504
rect 19852 16464 19858 16476
rect 5353 16439 5411 16445
rect 5353 16436 5365 16439
rect 4908 16408 5365 16436
rect 5353 16405 5365 16408
rect 5399 16436 5411 16439
rect 7006 16436 7012 16448
rect 5399 16408 7012 16436
rect 5399 16405 5411 16408
rect 5353 16399 5411 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 8415 16439 8473 16445
rect 8415 16405 8427 16439
rect 8461 16436 8473 16439
rect 9674 16436 9680 16448
rect 8461 16408 9680 16436
rect 8461 16405 8473 16408
rect 8415 16399 8473 16405
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 11422 16436 11428 16448
rect 9999 16408 11428 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16436 12127 16439
rect 13078 16436 13084 16448
rect 12115 16408 13084 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 17494 16396 17500 16448
rect 17552 16396 17558 16448
rect 19610 16396 19616 16448
rect 19668 16396 19674 16448
rect 19886 16396 19892 16448
rect 19944 16396 19950 16448
rect 19996 16436 20024 16476
rect 20990 16464 20996 16516
rect 21048 16464 21054 16516
rect 21174 16464 21180 16516
rect 21232 16464 21238 16516
rect 22020 16504 22048 16544
rect 22094 16532 22100 16584
rect 22152 16572 22158 16584
rect 22261 16575 22319 16581
rect 22261 16572 22273 16575
rect 22152 16544 22273 16572
rect 22152 16532 22158 16544
rect 22261 16541 22273 16544
rect 22307 16541 22319 16575
rect 23768 16572 23796 16680
rect 28258 16668 28264 16720
rect 28316 16668 28322 16720
rect 25130 16640 25136 16652
rect 24044 16612 25136 16640
rect 22261 16535 22319 16541
rect 23308 16544 23796 16572
rect 23308 16504 23336 16544
rect 23842 16532 23848 16584
rect 23900 16532 23906 16584
rect 24044 16581 24072 16612
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 26050 16640 26056 16652
rect 25240 16612 26056 16640
rect 24029 16575 24087 16581
rect 24029 16541 24041 16575
rect 24075 16541 24087 16575
rect 24029 16535 24087 16541
rect 24118 16532 24124 16584
rect 24176 16572 24182 16584
rect 24762 16572 24768 16584
rect 24176 16544 24768 16572
rect 24176 16532 24182 16544
rect 24762 16532 24768 16544
rect 24820 16532 24826 16584
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16572 24915 16575
rect 25240 16572 25268 16612
rect 26050 16600 26056 16612
rect 26108 16600 26114 16652
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 29104 16640 29132 16736
rect 29733 16643 29791 16649
rect 29733 16640 29745 16643
rect 26476 16612 27660 16640
rect 29104 16612 29745 16640
rect 26476 16600 26482 16612
rect 24903 16544 25268 16572
rect 27632 16572 27660 16612
rect 29733 16609 29745 16612
rect 29779 16609 29791 16643
rect 29733 16603 29791 16609
rect 28445 16575 28503 16581
rect 28445 16572 28457 16575
rect 27632 16544 28457 16572
rect 24903 16541 24915 16544
rect 24857 16535 24915 16541
rect 28445 16541 28457 16544
rect 28491 16541 28503 16575
rect 28445 16535 28503 16541
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 24136 16504 24164 16532
rect 22020 16476 23336 16504
rect 23400 16476 24164 16504
rect 25041 16507 25099 16513
rect 20070 16436 20076 16448
rect 19996 16408 20076 16436
rect 20070 16396 20076 16408
rect 20128 16436 20134 16448
rect 21192 16436 21220 16464
rect 22296 16448 22324 16476
rect 20128 16408 21220 16436
rect 20128 16396 20134 16408
rect 22278 16396 22284 16448
rect 22336 16396 22342 16448
rect 23400 16445 23428 16476
rect 25041 16473 25053 16507
rect 25087 16504 25099 16507
rect 25222 16504 25228 16516
rect 25087 16476 25228 16504
rect 25087 16473 25099 16476
rect 25041 16467 25099 16473
rect 25222 16464 25228 16476
rect 25280 16464 25286 16516
rect 26050 16464 26056 16516
rect 26108 16464 26114 16516
rect 28166 16464 28172 16516
rect 28224 16504 28230 16516
rect 28537 16507 28595 16513
rect 28537 16504 28549 16507
rect 28224 16476 28549 16504
rect 28224 16464 28230 16476
rect 28537 16473 28549 16476
rect 28583 16473 28595 16507
rect 28537 16467 28595 16473
rect 28626 16464 28632 16516
rect 28684 16464 28690 16516
rect 23385 16439 23443 16445
rect 23385 16405 23397 16439
rect 23431 16405 23443 16439
rect 23385 16399 23443 16405
rect 23934 16396 23940 16448
rect 23992 16396 23998 16448
rect 24394 16396 24400 16448
rect 24452 16436 24458 16448
rect 24581 16439 24639 16445
rect 24581 16436 24593 16439
rect 24452 16408 24593 16436
rect 24452 16396 24458 16408
rect 24581 16405 24593 16408
rect 24627 16405 24639 16439
rect 24581 16399 24639 16405
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 28828 16436 28856 16535
rect 29822 16532 29828 16584
rect 29880 16572 29886 16584
rect 29989 16575 30047 16581
rect 29989 16572 30001 16575
rect 29880 16544 30001 16572
rect 29880 16532 29886 16544
rect 29989 16541 30001 16544
rect 30035 16541 30047 16575
rect 29989 16535 30047 16541
rect 31846 16532 31852 16584
rect 31904 16532 31910 16584
rect 26292 16408 28856 16436
rect 26292 16396 26298 16408
rect 31662 16396 31668 16448
rect 31720 16396 31726 16448
rect 1104 16346 32632 16368
rect 1104 16294 8792 16346
rect 8844 16294 8856 16346
rect 8908 16294 8920 16346
rect 8972 16294 8984 16346
rect 9036 16294 9048 16346
rect 9100 16294 16634 16346
rect 16686 16294 16698 16346
rect 16750 16294 16762 16346
rect 16814 16294 16826 16346
rect 16878 16294 16890 16346
rect 16942 16294 24476 16346
rect 24528 16294 24540 16346
rect 24592 16294 24604 16346
rect 24656 16294 24668 16346
rect 24720 16294 24732 16346
rect 24784 16294 32318 16346
rect 32370 16294 32382 16346
rect 32434 16294 32446 16346
rect 32498 16294 32510 16346
rect 32562 16294 32574 16346
rect 32626 16294 32632 16346
rect 1104 16272 32632 16294
rect 1578 16192 1584 16244
rect 1636 16192 1642 16244
rect 2866 16192 2872 16244
rect 2924 16192 2930 16244
rect 3053 16235 3111 16241
rect 3053 16201 3065 16235
rect 3099 16232 3111 16235
rect 3099 16204 3924 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 2314 16124 2320 16176
rect 2372 16164 2378 16176
rect 3513 16167 3571 16173
rect 3513 16164 3525 16167
rect 2372 16136 3525 16164
rect 2372 16124 2378 16136
rect 3513 16133 3525 16136
rect 3559 16133 3571 16167
rect 3513 16127 3571 16133
rect 2038 16056 2044 16108
rect 2096 16096 2102 16108
rect 2501 16099 2559 16105
rect 2501 16096 2513 16099
rect 2096 16068 2513 16096
rect 2096 16056 2102 16068
rect 2501 16065 2513 16068
rect 2547 16096 2559 16099
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 2547 16068 3709 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 3786 16056 3792 16108
rect 3844 16056 3850 16108
rect 3896 16096 3924 16204
rect 4246 16192 4252 16244
rect 4304 16192 4310 16244
rect 5074 16192 5080 16244
rect 5132 16232 5138 16244
rect 8386 16232 8392 16244
rect 5132 16204 8392 16232
rect 5132 16192 5138 16204
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 5261 16167 5319 16173
rect 4120 16136 5212 16164
rect 4120 16124 4126 16136
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 3896 16068 4445 16096
rect 4433 16065 4445 16068
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16065 5043 16099
rect 5184 16096 5212 16136
rect 5261 16133 5273 16167
rect 5307 16164 5319 16167
rect 5721 16167 5779 16173
rect 5721 16164 5733 16167
rect 5307 16136 5733 16164
rect 5307 16133 5319 16136
rect 5261 16127 5319 16133
rect 5721 16133 5733 16136
rect 5767 16133 5779 16167
rect 6104 16164 6132 16204
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 10229 16235 10287 16241
rect 10229 16201 10241 16235
rect 10275 16232 10287 16235
rect 10962 16232 10968 16244
rect 10275 16204 10968 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 15197 16235 15255 16241
rect 15197 16232 15209 16235
rect 12584 16204 15209 16232
rect 12584 16192 12590 16204
rect 15197 16201 15209 16204
rect 15243 16201 15255 16235
rect 15197 16195 15255 16201
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 15712 16204 16865 16232
rect 15712 16192 15718 16204
rect 16853 16201 16865 16204
rect 16899 16201 16911 16235
rect 18627 16235 18685 16241
rect 18627 16232 18639 16235
rect 16853 16195 16911 16201
rect 18616 16201 18639 16232
rect 18673 16232 18685 16235
rect 19610 16232 19616 16244
rect 18673 16204 19616 16232
rect 18673 16201 18685 16204
rect 18616 16195 18685 16201
rect 7098 16164 7104 16176
rect 5721 16127 5779 16133
rect 6012 16136 6132 16164
rect 6656 16136 7104 16164
rect 6012 16105 6040 16136
rect 5997 16099 6055 16105
rect 5184 16068 5764 16096
rect 4985 16059 5043 16065
rect 3513 16031 3571 16037
rect 3513 15997 3525 16031
rect 3559 16028 3571 16031
rect 4062 16028 4068 16040
rect 3559 16000 4068 16028
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3528 15892 3556 15991
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 5000 16028 5028 16059
rect 5736 16037 5764 16068
rect 5997 16065 6009 16099
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 6656 16105 6684 16136
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 9582 16124 9588 16176
rect 9640 16124 9646 16176
rect 10318 16124 10324 16176
rect 10376 16164 10382 16176
rect 13354 16164 13360 16176
rect 10376 16136 13360 16164
rect 10376 16124 10382 16136
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 14642 16124 14648 16176
rect 14700 16124 14706 16176
rect 15565 16167 15623 16173
rect 15565 16133 15577 16167
rect 15611 16164 15623 16167
rect 16114 16164 16120 16176
rect 15611 16136 16120 16164
rect 15611 16133 15623 16136
rect 15565 16127 15623 16133
rect 16114 16124 16120 16136
rect 16172 16164 16178 16176
rect 16209 16167 16267 16173
rect 16209 16164 16221 16167
rect 16172 16136 16221 16164
rect 16172 16124 16178 16136
rect 16209 16133 16221 16136
rect 16255 16133 16267 16167
rect 16209 16127 16267 16133
rect 18414 16124 18420 16176
rect 18472 16124 18478 16176
rect 6641 16099 6699 16105
rect 6641 16096 6653 16099
rect 6144 16068 6653 16096
rect 6144 16056 6150 16068
rect 6641 16065 6653 16068
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 6730 16056 6736 16108
rect 6788 16056 6794 16108
rect 9214 16096 9220 16108
rect 6840 16068 9220 16096
rect 5721 16031 5779 16037
rect 5000 16000 5396 16028
rect 3602 15920 3608 15972
rect 3660 15960 3666 15972
rect 5074 15960 5080 15972
rect 3660 15932 5080 15960
rect 3660 15920 3666 15932
rect 5074 15920 5080 15932
rect 5132 15920 5138 15972
rect 5258 15920 5264 15972
rect 5316 15920 5322 15972
rect 5368 15960 5396 16000
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 6840 16028 6868 16068
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 11974 16096 11980 16108
rect 11808 16068 11980 16096
rect 5767 16000 6868 16028
rect 6917 16031 6975 16037
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 8294 16028 8300 16040
rect 6963 16000 8300 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 5905 15963 5963 15969
rect 5905 15960 5917 15963
rect 5368 15932 5917 15960
rect 5905 15929 5917 15932
rect 5951 15960 5963 15963
rect 6932 15960 6960 15991
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 8444 16000 11468 16028
rect 8444 15988 8450 16000
rect 5951 15932 6960 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 8536 15932 10057 15960
rect 8536 15920 8542 15932
rect 10045 15929 10057 15932
rect 10091 15929 10103 15963
rect 10045 15923 10103 15929
rect 10594 15920 10600 15972
rect 10652 15920 10658 15972
rect 11440 15960 11468 16000
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 11808 16028 11836 16068
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 13078 16096 13084 16108
rect 13035 16068 13084 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 13078 16056 13084 16068
rect 13136 16056 13142 16108
rect 13446 16056 13452 16108
rect 13504 16096 13510 16108
rect 15381 16099 15439 16105
rect 15381 16096 15393 16099
rect 13504 16068 15393 16096
rect 13504 16056 13510 16068
rect 15381 16065 15393 16068
rect 15427 16065 15439 16099
rect 15381 16059 15439 16065
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 15528 16068 15669 16096
rect 15528 16056 15534 16068
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 11572 16000 11836 16028
rect 11885 16031 11943 16037
rect 11572 15988 11578 16000
rect 11885 15997 11897 16031
rect 11931 16028 11943 16031
rect 12066 16028 12072 16040
rect 11931 16000 12072 16028
rect 11931 15997 11943 16000
rect 11885 15991 11943 15997
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 12158 15988 12164 16040
rect 12216 15988 12222 16040
rect 15838 16028 15844 16040
rect 13004 16000 15844 16028
rect 12176 15960 12204 15988
rect 13004 15972 13032 16000
rect 15838 15988 15844 16000
rect 15896 16028 15902 16040
rect 16316 16028 16344 16059
rect 17034 16056 17040 16108
rect 17092 16056 17098 16108
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 17770 16096 17776 16108
rect 17267 16068 17776 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 15896 16000 16344 16028
rect 17313 16031 17371 16037
rect 15896 15988 15902 16000
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 18616 16028 18644 16195
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 19702 16192 19708 16244
rect 19760 16192 19766 16244
rect 19978 16192 19984 16244
rect 20036 16232 20042 16244
rect 20073 16235 20131 16241
rect 20073 16232 20085 16235
rect 20036 16204 20085 16232
rect 20036 16192 20042 16204
rect 20073 16201 20085 16204
rect 20119 16201 20131 16235
rect 20073 16195 20131 16201
rect 20162 16192 20168 16244
rect 20220 16232 20226 16244
rect 23017 16235 23075 16241
rect 20220 16204 22094 16232
rect 20220 16192 20226 16204
rect 19889 16167 19947 16173
rect 19889 16133 19901 16167
rect 19935 16164 19947 16167
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 19935 16136 20821 16164
rect 19935 16133 19947 16136
rect 19889 16127 19947 16133
rect 20809 16133 20821 16136
rect 20855 16133 20867 16167
rect 22066 16164 22094 16204
rect 23017 16201 23029 16235
rect 23063 16232 23075 16235
rect 24026 16232 24032 16244
rect 23063 16204 24032 16232
rect 23063 16201 23075 16204
rect 23017 16195 23075 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 25409 16235 25467 16241
rect 25409 16201 25421 16235
rect 25455 16232 25467 16235
rect 25590 16232 25596 16244
rect 25455 16204 25596 16232
rect 25455 16201 25467 16204
rect 25409 16195 25467 16201
rect 25590 16192 25596 16204
rect 25648 16192 25654 16244
rect 27709 16235 27767 16241
rect 27709 16201 27721 16235
rect 27755 16232 27767 16235
rect 28626 16232 28632 16244
rect 27755 16204 28632 16232
rect 27755 16201 27767 16204
rect 27709 16195 27767 16201
rect 28626 16192 28632 16204
rect 28684 16192 28690 16244
rect 29730 16192 29736 16244
rect 29788 16192 29794 16244
rect 31757 16235 31815 16241
rect 31757 16201 31769 16235
rect 31803 16232 31815 16235
rect 31938 16232 31944 16244
rect 31803 16204 31944 16232
rect 31803 16201 31815 16204
rect 31757 16195 31815 16201
rect 31938 16192 31944 16204
rect 31996 16192 32002 16244
rect 22833 16167 22891 16173
rect 22066 16136 22784 16164
rect 20809 16127 20867 16133
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16096 20039 16099
rect 20070 16096 20076 16108
rect 20027 16068 20076 16096
rect 20027 16065 20039 16068
rect 19981 16059 20039 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 17359 16000 18644 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 20732 16028 20760 16059
rect 20898 16056 20904 16108
rect 20956 16056 20962 16108
rect 22756 16096 22784 16136
rect 22833 16133 22845 16167
rect 22879 16164 22891 16167
rect 23198 16164 23204 16176
rect 22879 16136 23204 16164
rect 22879 16133 22891 16136
rect 22833 16127 22891 16133
rect 23198 16124 23204 16136
rect 23256 16124 23262 16176
rect 23845 16167 23903 16173
rect 23845 16133 23857 16167
rect 23891 16164 23903 16167
rect 24118 16164 24124 16176
rect 23891 16136 24124 16164
rect 23891 16133 23903 16136
rect 23845 16127 23903 16133
rect 24118 16124 24124 16136
rect 24176 16124 24182 16176
rect 26602 16164 26608 16176
rect 24964 16136 26608 16164
rect 24964 16096 24992 16136
rect 22756 16068 24992 16096
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 25096 16068 25237 16096
rect 25096 16056 25102 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 25406 16056 25412 16108
rect 25464 16096 25470 16108
rect 26068 16105 26096 16136
rect 26602 16124 26608 16136
rect 26660 16124 26666 16176
rect 27614 16124 27620 16176
rect 27672 16164 27678 16176
rect 27672 16136 29224 16164
rect 27672 16124 27678 16136
rect 26053 16099 26111 16105
rect 25464 16068 26024 16096
rect 25464 16056 25470 16068
rect 21726 16028 21732 16040
rect 19944 16000 21732 16028
rect 19944 15988 19950 16000
rect 21726 15988 21732 16000
rect 21784 15988 21790 16040
rect 24949 16031 25007 16037
rect 24949 15997 24961 16031
rect 24995 15997 25007 16031
rect 24949 15991 25007 15997
rect 11440 15932 12204 15960
rect 12986 15920 12992 15972
rect 13044 15920 13050 15972
rect 18874 15920 18880 15972
rect 18932 15960 18938 15972
rect 18932 15932 19472 15960
rect 18932 15920 18938 15932
rect 2915 15864 3556 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 8110 15892 8116 15904
rect 7524 15864 8116 15892
rect 7524 15852 7530 15864
rect 8110 15852 8116 15864
rect 8168 15892 8174 15904
rect 8297 15895 8355 15901
rect 8297 15892 8309 15895
rect 8168 15864 8309 15892
rect 8168 15852 8174 15864
rect 8297 15861 8309 15864
rect 8343 15892 8355 15895
rect 9214 15892 9220 15904
rect 8343 15864 9220 15892
rect 8343 15861 8355 15864
rect 8297 15855 8355 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15892 10287 15895
rect 10502 15892 10508 15904
rect 10275 15864 10508 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 10502 15852 10508 15864
rect 10560 15892 10566 15904
rect 10686 15892 10692 15904
rect 10560 15864 10692 15892
rect 10560 15852 10566 15864
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11330 15852 11336 15904
rect 11388 15892 11394 15904
rect 11790 15892 11796 15904
rect 11388 15864 11796 15892
rect 11388 15852 11394 15864
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 12161 15895 12219 15901
rect 12161 15861 12173 15895
rect 12207 15892 12219 15895
rect 13170 15892 13176 15904
rect 12207 15864 13176 15892
rect 12207 15861 12219 15864
rect 12161 15855 12219 15861
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 18601 15895 18659 15901
rect 18601 15892 18613 15895
rect 16540 15864 18613 15892
rect 16540 15852 16546 15864
rect 18601 15861 18613 15864
rect 18647 15861 18659 15895
rect 18601 15855 18659 15861
rect 18785 15895 18843 15901
rect 18785 15861 18797 15895
rect 18831 15892 18843 15895
rect 19242 15892 19248 15904
rect 18831 15864 19248 15892
rect 18831 15861 18843 15864
rect 18785 15855 18843 15861
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 19444 15892 19472 15932
rect 19518 15920 19524 15972
rect 19576 15960 19582 15972
rect 20257 15963 20315 15969
rect 20257 15960 20269 15963
rect 19576 15932 20269 15960
rect 19576 15920 19582 15932
rect 20257 15929 20269 15932
rect 20303 15929 20315 15963
rect 22465 15963 22523 15969
rect 22465 15960 22477 15963
rect 20257 15923 20315 15929
rect 22066 15932 22477 15960
rect 20990 15892 20996 15904
rect 19444 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 21082 15852 21088 15904
rect 21140 15892 21146 15904
rect 22066 15892 22094 15932
rect 22465 15929 22477 15932
rect 22511 15929 22523 15963
rect 22465 15923 22523 15929
rect 23658 15920 23664 15972
rect 23716 15960 23722 15972
rect 24302 15960 24308 15972
rect 23716 15932 24308 15960
rect 23716 15920 23722 15932
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 24964 15904 24992 15991
rect 25866 15988 25872 16040
rect 25924 15988 25930 16040
rect 25996 16028 26024 16068
rect 26053 16065 26065 16099
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 26326 16056 26332 16108
rect 26384 16056 26390 16108
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16096 27399 16099
rect 28166 16096 28172 16108
rect 27387 16068 28172 16096
rect 27387 16065 27399 16068
rect 27341 16059 27399 16065
rect 27356 16028 27384 16059
rect 28166 16056 28172 16068
rect 28224 16056 28230 16108
rect 28276 16105 28304 16136
rect 28261 16099 28319 16105
rect 28261 16065 28273 16099
rect 28307 16065 28319 16099
rect 28261 16059 28319 16065
rect 28902 16056 28908 16108
rect 28960 16096 28966 16108
rect 29196 16105 29224 16136
rect 30374 16124 30380 16176
rect 30432 16164 30438 16176
rect 30432 16136 31616 16164
rect 30432 16124 30438 16136
rect 28997 16099 29055 16105
rect 28997 16096 29009 16099
rect 28960 16068 29009 16096
rect 28960 16056 28966 16068
rect 28997 16065 29009 16068
rect 29043 16065 29055 16099
rect 28997 16059 29055 16065
rect 29181 16099 29239 16105
rect 29181 16065 29193 16099
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 30857 16099 30915 16105
rect 30857 16065 30869 16099
rect 30903 16096 30915 16099
rect 31018 16096 31024 16108
rect 30903 16068 31024 16096
rect 30903 16065 30915 16068
rect 30857 16059 30915 16065
rect 31018 16056 31024 16068
rect 31076 16056 31082 16108
rect 31588 16105 31616 16136
rect 31573 16099 31631 16105
rect 31573 16065 31585 16099
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 25996 16000 27384 16028
rect 27433 16031 27491 16037
rect 27433 15997 27445 16031
rect 27479 16028 27491 16031
rect 29270 16028 29276 16040
rect 27479 16000 29276 16028
rect 27479 15997 27491 16000
rect 27433 15991 27491 15997
rect 25041 15963 25099 15969
rect 25041 15929 25053 15963
rect 25087 15960 25099 15963
rect 25130 15960 25136 15972
rect 25087 15932 25136 15960
rect 25087 15929 25099 15932
rect 25041 15923 25099 15929
rect 25130 15920 25136 15932
rect 25188 15960 25194 15972
rect 27448 15960 27476 15991
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 31110 15988 31116 16040
rect 31168 15988 31174 16040
rect 29089 15963 29147 15969
rect 29089 15960 29101 15963
rect 25188 15932 27476 15960
rect 27540 15932 29101 15960
rect 25188 15920 25194 15932
rect 21140 15864 22094 15892
rect 21140 15852 21146 15864
rect 22738 15852 22744 15904
rect 22796 15892 22802 15904
rect 22833 15895 22891 15901
rect 22833 15892 22845 15895
rect 22796 15864 22845 15892
rect 22796 15852 22802 15864
rect 22833 15861 22845 15864
rect 22879 15861 22891 15895
rect 22833 15855 22891 15861
rect 22922 15852 22928 15904
rect 22980 15892 22986 15904
rect 23569 15895 23627 15901
rect 23569 15892 23581 15895
rect 22980 15864 23581 15892
rect 22980 15852 22986 15864
rect 23569 15861 23581 15864
rect 23615 15861 23627 15895
rect 23569 15855 23627 15861
rect 24946 15852 24952 15904
rect 25004 15892 25010 15904
rect 27540 15892 27568 15932
rect 29089 15929 29101 15932
rect 29135 15929 29147 15963
rect 29089 15923 29147 15929
rect 25004 15864 27568 15892
rect 25004 15852 25010 15864
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 28445 15895 28503 15901
rect 28445 15892 28457 15895
rect 28224 15864 28457 15892
rect 28224 15852 28230 15864
rect 28445 15861 28457 15864
rect 28491 15861 28503 15895
rect 28445 15855 28503 15861
rect 1104 15802 32476 15824
rect 1104 15750 4871 15802
rect 4923 15750 4935 15802
rect 4987 15750 4999 15802
rect 5051 15750 5063 15802
rect 5115 15750 5127 15802
rect 5179 15750 12713 15802
rect 12765 15750 12777 15802
rect 12829 15750 12841 15802
rect 12893 15750 12905 15802
rect 12957 15750 12969 15802
rect 13021 15750 20555 15802
rect 20607 15750 20619 15802
rect 20671 15750 20683 15802
rect 20735 15750 20747 15802
rect 20799 15750 20811 15802
rect 20863 15750 28397 15802
rect 28449 15750 28461 15802
rect 28513 15750 28525 15802
rect 28577 15750 28589 15802
rect 28641 15750 28653 15802
rect 28705 15750 32476 15802
rect 1104 15728 32476 15750
rect 6086 15648 6092 15700
rect 6144 15648 6150 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8386 15688 8392 15700
rect 8067 15660 8392 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8628 15660 9321 15688
rect 8628 15648 8634 15660
rect 9309 15657 9321 15660
rect 9355 15688 9367 15691
rect 11238 15688 11244 15700
rect 9355 15660 11244 15688
rect 9355 15657 9367 15660
rect 9309 15651 9367 15657
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 11330 15648 11336 15700
rect 11388 15648 11394 15700
rect 11440 15660 14964 15688
rect 2866 15580 2872 15632
rect 2924 15620 2930 15632
rect 3602 15620 3608 15632
rect 2924 15592 3608 15620
rect 2924 15580 2930 15592
rect 3602 15580 3608 15592
rect 3660 15580 3666 15632
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 11440 15620 11468 15660
rect 10744 15592 11468 15620
rect 10744 15580 10750 15592
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 13173 15623 13231 15629
rect 13173 15620 13185 15623
rect 11664 15592 13185 15620
rect 11664 15580 11670 15592
rect 13173 15589 13185 15592
rect 13219 15620 13231 15623
rect 14366 15620 14372 15632
rect 13219 15592 14372 15620
rect 13219 15589 13231 15592
rect 13173 15583 13231 15589
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 14936 15620 14964 15660
rect 15102 15648 15108 15700
rect 15160 15648 15166 15700
rect 15933 15691 15991 15697
rect 15933 15657 15945 15691
rect 15979 15688 15991 15691
rect 16482 15688 16488 15700
rect 15979 15660 16488 15688
rect 15979 15657 15991 15660
rect 15933 15651 15991 15657
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 17037 15691 17095 15697
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 17678 15688 17684 15700
rect 17083 15660 17684 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 17773 15691 17831 15697
rect 17773 15657 17785 15691
rect 17819 15688 17831 15691
rect 18506 15688 18512 15700
rect 17819 15660 18512 15688
rect 17819 15657 17831 15660
rect 17773 15651 17831 15657
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 19610 15688 19616 15700
rect 18739 15660 19616 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 21082 15648 21088 15700
rect 21140 15648 21146 15700
rect 21177 15691 21235 15697
rect 21177 15657 21189 15691
rect 21223 15688 21235 15691
rect 21358 15688 21364 15700
rect 21223 15660 21364 15688
rect 21223 15657 21235 15660
rect 21177 15651 21235 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21818 15648 21824 15700
rect 21876 15648 21882 15700
rect 23198 15648 23204 15700
rect 23256 15648 23262 15700
rect 25038 15648 25044 15700
rect 25096 15648 25102 15700
rect 25314 15648 25320 15700
rect 25372 15688 25378 15700
rect 25372 15660 25544 15688
rect 25372 15648 25378 15660
rect 18877 15623 18935 15629
rect 14936 15592 18000 15620
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15552 2743 15555
rect 4062 15552 4068 15564
rect 2731 15524 4068 15552
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 7466 15512 7472 15564
rect 7524 15512 7530 15564
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11514 15552 11520 15564
rect 11296 15524 11520 15552
rect 11296 15512 11302 15524
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 12618 15552 12624 15564
rect 12575 15524 12624 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 13771 15524 16896 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 3234 15484 3240 15496
rect 2639 15456 3240 15484
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15484 3479 15487
rect 3786 15484 3792 15496
rect 3467 15456 3792 15484
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 8202 15444 8208 15496
rect 8260 15444 8266 15496
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10689 15487 10747 15493
rect 10192 15456 10548 15484
rect 10192 15444 10198 15456
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15416 1823 15419
rect 3510 15416 3516 15428
rect 1811 15388 3516 15416
rect 1811 15385 1823 15388
rect 1765 15379 1823 15385
rect 3510 15376 3516 15388
rect 3568 15376 3574 15428
rect 7224 15419 7282 15425
rect 7224 15385 7236 15419
rect 7270 15416 7282 15419
rect 8386 15416 8392 15428
rect 7270 15388 8392 15416
rect 7270 15385 7282 15388
rect 7224 15379 7282 15385
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 8570 15376 8576 15428
rect 8628 15416 8634 15428
rect 10422 15419 10480 15425
rect 10422 15416 10434 15419
rect 8628 15388 10434 15416
rect 8628 15376 8634 15388
rect 10422 15385 10434 15388
rect 10468 15385 10480 15419
rect 10520 15416 10548 15456
rect 10689 15453 10701 15487
rect 10735 15484 10747 15487
rect 11882 15484 11888 15496
rect 10735 15456 11888 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 12158 15444 12164 15496
rect 12216 15444 12222 15496
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12308 15456 12357 15484
rect 12308 15444 12314 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15484 12771 15487
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 12759 15456 13461 15484
rect 12759 15453 12771 15456
rect 12713 15447 12771 15453
rect 13449 15453 13461 15456
rect 13495 15484 13507 15487
rect 13630 15484 13636 15496
rect 13495 15456 13636 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 13630 15444 13636 15456
rect 13688 15484 13694 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 13688 15456 14841 15484
rect 13688 15444 13694 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 15252 15456 15577 15484
rect 15252 15444 15258 15456
rect 15565 15453 15577 15456
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 16868 15493 16896 15524
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 17972 15484 18000 15592
rect 18877 15589 18889 15623
rect 18923 15620 18935 15623
rect 21100 15620 21128 15648
rect 18923 15592 21128 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 18892 15552 18920 15583
rect 21726 15580 21732 15632
rect 21784 15620 21790 15632
rect 25516 15620 25544 15660
rect 27430 15648 27436 15700
rect 27488 15688 27494 15700
rect 28534 15688 28540 15700
rect 27488 15660 28540 15688
rect 27488 15648 27494 15660
rect 28534 15648 28540 15660
rect 28592 15688 28598 15700
rect 28629 15691 28687 15697
rect 28629 15688 28641 15691
rect 28592 15660 28641 15688
rect 28592 15648 28598 15660
rect 28629 15657 28641 15660
rect 28675 15657 28687 15691
rect 28629 15651 28687 15657
rect 28736 15660 28994 15688
rect 25774 15620 25780 15632
rect 21784 15592 23152 15620
rect 21784 15580 21790 15592
rect 18748 15524 18920 15552
rect 18748 15512 18754 15524
rect 19150 15512 19156 15564
rect 19208 15552 19214 15564
rect 20162 15552 20168 15564
rect 19208 15524 20168 15552
rect 19208 15512 19214 15524
rect 17972 15456 19196 15484
rect 11301 15419 11359 15425
rect 11301 15416 11313 15419
rect 10520 15388 11313 15416
rect 10422 15379 10480 15385
rect 11301 15385 11313 15388
rect 11347 15385 11359 15419
rect 11301 15379 11359 15385
rect 11514 15376 11520 15428
rect 11572 15376 11578 15428
rect 13354 15376 13360 15428
rect 13412 15416 13418 15428
rect 13906 15416 13912 15428
rect 13412 15388 13912 15416
rect 13412 15376 13418 15388
rect 13906 15376 13912 15388
rect 13964 15416 13970 15428
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 13964 15388 14381 15416
rect 13964 15376 13970 15388
rect 14369 15385 14381 15388
rect 14415 15416 14427 15419
rect 14458 15416 14464 15428
rect 14415 15388 14464 15416
rect 14415 15385 14427 15388
rect 14369 15379 14427 15385
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 17972 15425 18000 15456
rect 14921 15419 14979 15425
rect 14921 15385 14933 15419
rect 14967 15416 14979 15419
rect 17957 15419 18015 15425
rect 14967 15388 17908 15416
rect 14967 15385 14979 15388
rect 14921 15379 14979 15385
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 2225 15351 2283 15357
rect 2225 15348 2237 15351
rect 2188 15320 2237 15348
rect 2188 15308 2194 15320
rect 2225 15317 2237 15320
rect 2271 15317 2283 15351
rect 2225 15311 2283 15317
rect 3329 15351 3387 15357
rect 3329 15317 3341 15351
rect 3375 15348 3387 15351
rect 3602 15348 3608 15360
rect 3375 15320 3608 15348
rect 3375 15317 3387 15320
rect 3329 15311 3387 15317
rect 3602 15308 3608 15320
rect 3660 15308 3666 15360
rect 10594 15308 10600 15360
rect 10652 15348 10658 15360
rect 11149 15351 11207 15357
rect 11149 15348 11161 15351
rect 10652 15320 11161 15348
rect 10652 15308 10658 15320
rect 11149 15317 11161 15320
rect 11195 15317 11207 15351
rect 11149 15311 11207 15317
rect 13538 15308 13544 15360
rect 13596 15308 13602 15360
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 16482 15348 16488 15360
rect 15528 15320 16488 15348
rect 15528 15308 15534 15320
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 17770 15357 17776 15360
rect 17589 15351 17647 15357
rect 17589 15348 17601 15351
rect 17368 15320 17601 15348
rect 17368 15308 17374 15320
rect 17589 15317 17601 15320
rect 17635 15317 17647 15351
rect 17589 15311 17647 15317
rect 17757 15351 17776 15357
rect 17757 15317 17769 15351
rect 17757 15311 17776 15317
rect 17770 15308 17776 15311
rect 17828 15308 17834 15360
rect 17880 15348 17908 15388
rect 17957 15385 17969 15419
rect 18003 15385 18015 15419
rect 17957 15379 18015 15385
rect 18414 15376 18420 15428
rect 18472 15416 18478 15428
rect 18509 15419 18567 15425
rect 18509 15416 18521 15419
rect 18472 15388 18521 15416
rect 18472 15376 18478 15388
rect 18509 15385 18521 15388
rect 18555 15385 18567 15419
rect 19168 15416 19196 15456
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 19536 15493 19564 15524
rect 20162 15512 20168 15524
rect 20220 15512 20226 15564
rect 20898 15552 20904 15564
rect 20364 15524 20904 15552
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19300 15456 19441 15484
rect 19300 15444 19306 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19668 15456 19717 15484
rect 19668 15444 19674 15456
rect 19705 15453 19717 15456
rect 19751 15484 19763 15487
rect 20364 15484 20392 15524
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 22922 15552 22928 15564
rect 21376 15524 22928 15552
rect 19751 15456 20392 15484
rect 19751 15453 19763 15456
rect 19705 15447 19763 15453
rect 20438 15444 20444 15496
rect 20496 15484 20502 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20496 15456 20545 15484
rect 20496 15444 20502 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 21376 15484 21404 15524
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 21048 15456 21404 15484
rect 21048 15444 21054 15456
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21692 15456 22017 15484
rect 21692 15444 21698 15456
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 22005 15447 22063 15453
rect 22189 15487 22247 15493
rect 22189 15453 22201 15487
rect 22235 15484 22247 15487
rect 22278 15484 22284 15496
rect 22235 15456 22284 15484
rect 22235 15453 22247 15456
rect 22189 15447 22247 15453
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 23124 15484 23152 15592
rect 23400 15592 23888 15620
rect 25516 15592 25780 15620
rect 23198 15512 23204 15564
rect 23256 15552 23262 15564
rect 23400 15561 23428 15592
rect 23385 15555 23443 15561
rect 23385 15552 23397 15555
rect 23256 15524 23397 15552
rect 23256 15512 23262 15524
rect 23385 15521 23397 15524
rect 23431 15521 23443 15555
rect 23658 15552 23664 15564
rect 23620 15524 23664 15552
rect 23385 15515 23443 15521
rect 23658 15512 23664 15524
rect 23716 15512 23722 15564
rect 23860 15552 23888 15592
rect 25774 15580 25780 15592
rect 25832 15620 25838 15632
rect 26786 15620 26792 15632
rect 25832 15592 26792 15620
rect 25832 15580 25838 15592
rect 26786 15580 26792 15592
rect 26844 15620 26850 15632
rect 28736 15620 28764 15660
rect 26844 15592 28764 15620
rect 28813 15623 28871 15629
rect 26844 15580 26850 15592
rect 28813 15589 28825 15623
rect 28859 15589 28871 15623
rect 28966 15620 28994 15660
rect 29270 15648 29276 15700
rect 29328 15688 29334 15700
rect 30469 15691 30527 15697
rect 30469 15688 30481 15691
rect 29328 15660 30481 15688
rect 29328 15648 29334 15660
rect 30469 15657 30481 15660
rect 30515 15657 30527 15691
rect 30469 15651 30527 15657
rect 31018 15648 31024 15700
rect 31076 15648 31082 15700
rect 28966 15592 30328 15620
rect 28813 15583 28871 15589
rect 23934 15552 23940 15564
rect 23860 15524 23940 15552
rect 23934 15512 23940 15524
rect 23992 15552 23998 15564
rect 28261 15555 28319 15561
rect 28261 15552 28273 15555
rect 23992 15524 28273 15552
rect 23992 15512 23998 15524
rect 28261 15521 28273 15524
rect 28307 15521 28319 15555
rect 28828 15552 28856 15583
rect 30190 15552 30196 15564
rect 28828 15524 30196 15552
rect 28261 15515 28319 15521
rect 30190 15512 30196 15524
rect 30248 15512 30254 15564
rect 30300 15500 30328 15592
rect 30374 15580 30380 15632
rect 30432 15620 30438 15632
rect 30432 15592 31248 15620
rect 30432 15580 30438 15592
rect 30377 15500 30435 15503
rect 30300 15497 30435 15500
rect 23474 15484 23480 15496
rect 23124 15456 23480 15484
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 23750 15484 23756 15496
rect 23615 15456 23756 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 23750 15444 23756 15456
rect 23808 15484 23814 15496
rect 23808 15456 25176 15484
rect 23808 15444 23814 15456
rect 20806 15416 20812 15428
rect 19168 15388 20812 15416
rect 18509 15379 18567 15385
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 21726 15376 21732 15428
rect 21784 15376 21790 15428
rect 22738 15416 22744 15428
rect 22296 15388 22744 15416
rect 18322 15348 18328 15360
rect 17880 15320 18328 15348
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 18598 15308 18604 15360
rect 18656 15348 18662 15360
rect 18719 15351 18777 15357
rect 18719 15348 18731 15351
rect 18656 15320 18731 15348
rect 18656 15308 18662 15320
rect 18719 15317 18731 15320
rect 18765 15348 18777 15351
rect 19150 15348 19156 15360
rect 18765 15320 19156 15348
rect 18765 15317 18777 15320
rect 18719 15311 18777 15317
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 20254 15348 20260 15360
rect 19935 15320 20260 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 20346 15308 20352 15360
rect 20404 15308 20410 15360
rect 20824 15348 20852 15376
rect 22296 15348 22324 15388
rect 22738 15376 22744 15388
rect 22796 15416 22802 15428
rect 24854 15416 24860 15428
rect 22796 15388 24860 15416
rect 22796 15376 22802 15388
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 25148 15416 25176 15456
rect 25222 15444 25228 15496
rect 25280 15444 25286 15496
rect 25314 15444 25320 15496
rect 25372 15444 25378 15496
rect 25406 15444 25412 15496
rect 25464 15444 25470 15496
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15484 25559 15487
rect 25682 15484 25688 15496
rect 25547 15456 25688 15484
rect 25547 15453 25559 15456
rect 25501 15447 25559 15453
rect 25516 15416 25544 15447
rect 25682 15444 25688 15456
rect 25740 15444 25746 15496
rect 26050 15444 26056 15496
rect 26108 15444 26114 15496
rect 28994 15444 29000 15496
rect 29052 15484 29058 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29052 15456 29745 15484
rect 29052 15444 29058 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15484 29975 15487
rect 30006 15484 30012 15496
rect 29963 15456 30012 15484
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 30006 15444 30012 15456
rect 30064 15444 30070 15496
rect 30300 15472 30389 15497
rect 30377 15463 30389 15472
rect 30423 15463 30435 15497
rect 31220 15493 31248 15592
rect 30377 15457 30435 15463
rect 30561 15487 30619 15493
rect 30561 15453 30573 15487
rect 30607 15453 30619 15487
rect 30561 15447 30619 15453
rect 31205 15487 31263 15493
rect 31205 15453 31217 15487
rect 31251 15453 31263 15487
rect 31205 15447 31263 15453
rect 25148 15388 25544 15416
rect 28629 15419 28687 15425
rect 28629 15385 28641 15419
rect 28675 15416 28687 15419
rect 29825 15419 29883 15425
rect 29825 15416 29837 15419
rect 28675 15388 29837 15416
rect 28675 15385 28687 15388
rect 28629 15379 28687 15385
rect 29825 15385 29837 15388
rect 29871 15385 29883 15419
rect 29825 15379 29883 15385
rect 30098 15376 30104 15428
rect 30156 15416 30162 15428
rect 30576 15416 30604 15447
rect 30156 15388 30604 15416
rect 30156 15376 30162 15388
rect 20824 15320 22324 15348
rect 22373 15351 22431 15357
rect 22373 15317 22385 15351
rect 22419 15348 22431 15351
rect 24302 15348 24308 15360
rect 22419 15320 24308 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 24302 15308 24308 15320
rect 24360 15308 24366 15360
rect 24872 15348 24900 15376
rect 27430 15348 27436 15360
rect 24872 15320 27436 15348
rect 27430 15308 27436 15320
rect 27488 15308 27494 15360
rect 27525 15351 27583 15357
rect 27525 15317 27537 15351
rect 27571 15348 27583 15351
rect 27706 15348 27712 15360
rect 27571 15320 27712 15348
rect 27571 15317 27583 15320
rect 27525 15311 27583 15317
rect 27706 15308 27712 15320
rect 27764 15308 27770 15360
rect 28534 15308 28540 15360
rect 28592 15348 28598 15360
rect 30374 15348 30380 15360
rect 28592 15320 30380 15348
rect 28592 15308 28598 15320
rect 30374 15308 30380 15320
rect 30432 15348 30438 15360
rect 31662 15348 31668 15360
rect 30432 15320 31668 15348
rect 30432 15308 30438 15320
rect 31662 15308 31668 15320
rect 31720 15308 31726 15360
rect 1104 15258 32632 15280
rect 1104 15206 8792 15258
rect 8844 15206 8856 15258
rect 8908 15206 8920 15258
rect 8972 15206 8984 15258
rect 9036 15206 9048 15258
rect 9100 15206 16634 15258
rect 16686 15206 16698 15258
rect 16750 15206 16762 15258
rect 16814 15206 16826 15258
rect 16878 15206 16890 15258
rect 16942 15206 24476 15258
rect 24528 15206 24540 15258
rect 24592 15206 24604 15258
rect 24656 15206 24668 15258
rect 24720 15206 24732 15258
rect 24784 15206 32318 15258
rect 32370 15206 32382 15258
rect 32434 15206 32446 15258
rect 32498 15206 32510 15258
rect 32562 15206 32574 15258
rect 32626 15206 32632 15258
rect 1104 15184 32632 15206
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8570 15144 8576 15156
rect 8251 15116 8576 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 16114 15104 16120 15156
rect 16172 15104 16178 15156
rect 17037 15147 17095 15153
rect 17037 15144 17049 15147
rect 16224 15116 17049 15144
rect 8941 15079 8999 15085
rect 8941 15045 8953 15079
rect 8987 15076 8999 15079
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 8987 15048 9413 15076
rect 8987 15045 8999 15048
rect 8941 15039 8999 15045
rect 9401 15045 9413 15048
rect 9447 15045 9459 15079
rect 9401 15039 9459 15045
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10505 15079 10563 15085
rect 10505 15076 10517 15079
rect 10008 15048 10517 15076
rect 10008 15036 10014 15048
rect 10505 15045 10517 15048
rect 10551 15045 10563 15079
rect 10505 15039 10563 15045
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11974 15076 11980 15088
rect 11480 15048 11980 15076
rect 11480 15036 11486 15048
rect 11974 15036 11980 15048
rect 12032 15076 12038 15088
rect 12032 15048 15332 15076
rect 12032 15036 12038 15048
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 15008 2559 15011
rect 3050 15008 3056 15020
rect 2547 14980 3056 15008
rect 2547 14977 2559 14980
rect 2501 14971 2559 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 15008 3571 15011
rect 3970 15008 3976 15020
rect 3559 14980 3976 15008
rect 3559 14977 3571 14980
rect 3513 14971 3571 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7098 15008 7104 15020
rect 6963 14980 7104 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8478 15008 8484 15020
rect 8067 14980 8484 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8662 14968 8668 15020
rect 8720 14968 8726 15020
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 15008 8815 15011
rect 9674 15008 9680 15020
rect 8803 14980 9680 15008
rect 8803 14977 8815 14980
rect 8757 14971 8815 14977
rect 9674 14968 9680 14980
rect 9732 15008 9738 15020
rect 11698 15008 11704 15020
rect 9732 14980 11704 15008
rect 9732 14968 9738 14980
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 12492 14980 13185 15008
rect 12492 14968 12498 14980
rect 13173 14977 13185 14980
rect 13219 15008 13231 15011
rect 13538 15008 13544 15020
rect 13219 14980 13544 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 13630 14968 13636 15020
rect 13688 14968 13694 15020
rect 13906 14968 13912 15020
rect 13964 14968 13970 15020
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14424 14980 14473 15008
rect 14424 14968 14430 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 15102 14968 15108 15020
rect 15160 14968 15166 15020
rect 15304 15017 15332 15048
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15378 14968 15384 15020
rect 15436 14968 15442 15020
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16224 15008 16252 15116
rect 17037 15113 17049 15116
rect 17083 15144 17095 15147
rect 17770 15144 17776 15156
rect 17083 15116 17776 15144
rect 17083 15113 17095 15116
rect 17037 15107 17095 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18506 15104 18512 15156
rect 18564 15104 18570 15156
rect 22186 15144 22192 15156
rect 18616 15116 22192 15144
rect 16301 15079 16359 15085
rect 16301 15045 16313 15079
rect 16347 15076 16359 15079
rect 17589 15079 17647 15085
rect 17589 15076 17601 15079
rect 16347 15048 17601 15076
rect 16347 15045 16359 15048
rect 16301 15039 16359 15045
rect 17589 15045 17601 15048
rect 17635 15045 17647 15079
rect 18616 15076 18644 15116
rect 22186 15104 22192 15116
rect 22244 15144 22250 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 22244 15116 22293 15144
rect 22244 15104 22250 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22281 15107 22339 15113
rect 23124 15116 24164 15144
rect 17589 15039 17647 15045
rect 17696 15048 18644 15076
rect 19521 15079 19579 15085
rect 16071 14980 16252 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16540 14980 16865 15008
rect 16540 14968 16546 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17696 15008 17724 15048
rect 19521 15045 19533 15079
rect 19567 15076 19579 15079
rect 20593 15079 20651 15085
rect 20593 15076 20605 15079
rect 19567 15048 20605 15076
rect 19567 15045 19579 15048
rect 19521 15039 19579 15045
rect 20593 15045 20605 15048
rect 20639 15045 20651 15079
rect 20593 15039 20651 15045
rect 20806 15036 20812 15088
rect 20864 15036 20870 15088
rect 21450 15036 21456 15088
rect 21508 15076 21514 15088
rect 21508 15048 22508 15076
rect 21508 15036 21514 15048
rect 17175 14980 17724 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 2590 14900 2596 14952
rect 2648 14900 2654 14952
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 6086 14940 6092 14952
rect 3651 14912 6092 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 6086 14900 6092 14912
rect 6144 14940 6150 14952
rect 6638 14940 6644 14952
rect 6144 14912 6644 14940
rect 6144 14900 6150 14912
rect 6638 14900 6644 14912
rect 6696 14900 6702 14952
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 7239 14912 9413 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 9401 14909 9413 14912
rect 9447 14940 9459 14943
rect 13354 14940 13360 14952
rect 9447 14912 13360 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 13354 14900 13360 14912
rect 13412 14940 13418 14952
rect 13722 14940 13728 14952
rect 13412 14912 13728 14940
rect 13412 14900 13418 14912
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 14090 14900 14096 14952
rect 14148 14900 14154 14952
rect 17144 14940 17172 14971
rect 17770 14968 17776 15020
rect 17828 14968 17834 15020
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 15008 18107 15011
rect 19242 15008 19248 15020
rect 18095 14980 19248 15008
rect 18095 14977 18107 14980
rect 18049 14971 18107 14977
rect 19242 14968 19248 14980
rect 19300 15008 19306 15020
rect 19889 15011 19947 15017
rect 19889 15008 19901 15011
rect 19300 14980 19901 15008
rect 19300 14968 19306 14980
rect 19889 14977 19901 14980
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20162 15008 20168 15020
rect 20027 14980 20168 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20438 14968 20444 15020
rect 20496 14968 20502 15020
rect 22370 14968 22376 15020
rect 22428 14968 22434 15020
rect 22480 15017 22508 15048
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 15008 22891 15011
rect 23124 15008 23152 15116
rect 23566 15036 23572 15088
rect 23624 15076 23630 15088
rect 24136 15085 24164 15116
rect 24210 15104 24216 15156
rect 24268 15144 24274 15156
rect 24673 15147 24731 15153
rect 24673 15144 24685 15147
rect 24268 15116 24685 15144
rect 24268 15104 24274 15116
rect 24673 15113 24685 15116
rect 24719 15113 24731 15147
rect 24673 15107 24731 15113
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 26234 15104 26240 15156
rect 26292 15144 26298 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 26292 15116 27169 15144
rect 26292 15104 26298 15116
rect 27157 15113 27169 15116
rect 27203 15113 27215 15147
rect 27157 15107 27215 15113
rect 28353 15147 28411 15153
rect 28353 15113 28365 15147
rect 28399 15144 28411 15147
rect 28718 15144 28724 15156
rect 28399 15116 28724 15144
rect 28399 15113 28411 15116
rect 28353 15107 28411 15113
rect 28718 15104 28724 15116
rect 28776 15104 28782 15156
rect 29457 15147 29515 15153
rect 29457 15113 29469 15147
rect 29503 15144 29515 15147
rect 29730 15144 29736 15156
rect 29503 15116 29736 15144
rect 29503 15113 29515 15116
rect 29457 15107 29515 15113
rect 29730 15104 29736 15116
rect 29788 15104 29794 15156
rect 24121 15079 24179 15085
rect 23624 15048 23980 15076
rect 23624 15036 23630 15048
rect 22879 14980 23152 15008
rect 22879 14977 22891 14980
rect 22833 14971 22891 14977
rect 23198 14968 23204 15020
rect 23256 14968 23262 15020
rect 23290 14968 23296 15020
rect 23348 15008 23354 15020
rect 23952 15017 23980 15048
rect 24121 15045 24133 15079
rect 24167 15076 24179 15079
rect 24964 15076 24992 15104
rect 24167 15048 24992 15076
rect 24167 15045 24179 15048
rect 24121 15039 24179 15045
rect 25130 15036 25136 15088
rect 25188 15076 25194 15088
rect 27309 15079 27367 15085
rect 27309 15076 27321 15079
rect 25188 15048 27321 15076
rect 25188 15036 25194 15048
rect 27309 15045 27321 15048
rect 27355 15045 27367 15079
rect 27309 15039 27367 15045
rect 27430 15036 27436 15088
rect 27488 15076 27494 15088
rect 27525 15079 27583 15085
rect 27525 15076 27537 15079
rect 27488 15048 27537 15076
rect 27488 15036 27494 15048
rect 27525 15045 27537 15048
rect 27571 15045 27583 15079
rect 27525 15039 27583 15045
rect 27985 15079 28043 15085
rect 27985 15045 27997 15079
rect 28031 15076 28043 15079
rect 28074 15076 28080 15088
rect 28031 15048 28080 15076
rect 28031 15045 28043 15048
rect 27985 15039 28043 15045
rect 28074 15036 28080 15048
rect 28132 15036 28138 15088
rect 28258 15085 28264 15088
rect 28201 15079 28264 15085
rect 28201 15045 28213 15079
rect 28247 15045 28264 15079
rect 28201 15039 28264 15045
rect 28258 15036 28264 15039
rect 28316 15076 28322 15088
rect 30006 15076 30012 15088
rect 28316 15048 30012 15076
rect 28316 15036 28322 15048
rect 30006 15036 30012 15048
rect 30064 15036 30070 15088
rect 31110 15036 31116 15088
rect 31168 15076 31174 15088
rect 31168 15048 31708 15076
rect 31168 15036 31174 15048
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23348 14980 23857 15008
rect 23348 14968 23354 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 24854 14968 24860 15020
rect 24912 15008 24918 15020
rect 24949 15011 25007 15017
rect 24949 15008 24961 15011
rect 24912 14980 24961 15008
rect 24912 14968 24918 14980
rect 24949 14977 24961 14980
rect 24995 14977 25007 15011
rect 24949 14971 25007 14977
rect 25774 14968 25780 15020
rect 25832 14968 25838 15020
rect 25958 14968 25964 15020
rect 26016 15008 26022 15020
rect 26053 15011 26111 15017
rect 26053 15008 26065 15011
rect 26016 14980 26065 15008
rect 26016 14968 26022 14980
rect 26053 14977 26065 14980
rect 26099 15008 26111 15011
rect 26326 15008 26332 15020
rect 26099 14980 26332 15008
rect 26099 14977 26111 14980
rect 26053 14971 26111 14977
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 26510 14968 26516 15020
rect 26568 15008 26574 15020
rect 26568 14980 29040 15008
rect 26568 14968 26574 14980
rect 14752 14912 17172 14940
rect 17972 14940 18000 14968
rect 18598 14940 18604 14952
rect 17972 14912 18604 14940
rect 2869 14875 2927 14881
rect 2869 14841 2881 14875
rect 2915 14872 2927 14875
rect 5626 14872 5632 14884
rect 2915 14844 5632 14872
rect 2915 14841 2927 14844
rect 2869 14835 2927 14841
rect 5626 14832 5632 14844
rect 5684 14832 5690 14884
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7009 14875 7067 14881
rect 7009 14872 7021 14875
rect 6972 14844 7021 14872
rect 6972 14832 6978 14844
rect 7009 14841 7021 14844
rect 7055 14841 7067 14875
rect 7009 14835 7067 14841
rect 10134 14832 10140 14884
rect 10192 14832 10198 14884
rect 11882 14832 11888 14884
rect 11940 14872 11946 14884
rect 14642 14872 14648 14884
rect 11940 14844 14648 14872
rect 11940 14832 11946 14844
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 4522 14804 4528 14816
rect 3835 14776 4528 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 7101 14807 7159 14813
rect 7101 14773 7113 14807
rect 7147 14804 7159 14807
rect 8110 14804 8116 14816
rect 7147 14776 8116 14804
rect 7147 14773 7159 14776
rect 7101 14767 7159 14773
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 8941 14807 8999 14813
rect 8941 14773 8953 14807
rect 8987 14804 8999 14807
rect 9306 14804 9312 14816
rect 8987 14776 9312 14804
rect 8987 14773 8999 14776
rect 8941 14767 8999 14773
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 9582 14764 9588 14816
rect 9640 14764 9646 14816
rect 10502 14764 10508 14816
rect 10560 14764 10566 14816
rect 10686 14764 10692 14816
rect 10744 14764 10750 14816
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 14752 14804 14780 14912
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 18782 14900 18788 14952
rect 18840 14900 18846 14952
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 15746 14872 15752 14884
rect 15396 14844 15752 14872
rect 15396 14813 15424 14844
rect 15746 14832 15752 14844
rect 15804 14832 15810 14884
rect 17034 14872 17040 14884
rect 16224 14844 17040 14872
rect 13688 14776 14780 14804
rect 15381 14807 15439 14813
rect 13688 14764 13694 14776
rect 15381 14773 15393 14807
rect 15427 14773 15439 14807
rect 15381 14767 15439 14773
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14804 15623 14807
rect 16224 14804 16252 14844
rect 17034 14832 17040 14844
rect 17092 14832 17098 14884
rect 18892 14872 18920 14903
rect 18966 14900 18972 14952
rect 19024 14900 19030 14952
rect 19150 14900 19156 14952
rect 19208 14940 19214 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19208 14912 19625 14940
rect 19208 14900 19214 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 19702 14900 19708 14952
rect 19760 14900 19766 14952
rect 19978 14872 19984 14884
rect 18892 14844 19984 14872
rect 15611 14776 16252 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 16298 14764 16304 14816
rect 16356 14764 16362 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17126 14804 17132 14816
rect 17000 14776 17132 14804
rect 17000 14764 17006 14776
rect 17126 14764 17132 14776
rect 17184 14804 17190 14816
rect 18892 14804 18920 14844
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 20456 14881 20484 14968
rect 21634 14900 21640 14952
rect 21692 14940 21698 14952
rect 25685 14943 25743 14949
rect 21692 14912 23796 14940
rect 21692 14900 21698 14912
rect 20441 14875 20499 14881
rect 20441 14841 20453 14875
rect 20487 14841 20499 14875
rect 20441 14835 20499 14841
rect 17184 14776 18920 14804
rect 17184 14764 17190 14776
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 20312 14776 20637 14804
rect 20312 14764 20318 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 20625 14767 20683 14773
rect 22462 14764 22468 14816
rect 22520 14804 22526 14816
rect 23661 14807 23719 14813
rect 23661 14804 23673 14807
rect 22520 14776 23673 14804
rect 22520 14764 22526 14776
rect 23661 14773 23673 14776
rect 23707 14773 23719 14807
rect 23768 14804 23796 14912
rect 25685 14909 25697 14943
rect 25731 14940 25743 14943
rect 25866 14940 25872 14952
rect 25731 14912 25872 14940
rect 25731 14909 25743 14912
rect 25685 14903 25743 14909
rect 25866 14900 25872 14912
rect 25924 14900 25930 14952
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14940 26203 14943
rect 28902 14940 28908 14952
rect 26191 14912 28908 14940
rect 26191 14909 26203 14912
rect 26145 14903 26203 14909
rect 28902 14900 28908 14912
rect 28960 14900 28966 14952
rect 29012 14940 29040 14980
rect 29362 14968 29368 15020
rect 29420 14968 29426 15020
rect 30466 15008 30472 15020
rect 29472 14980 30472 15008
rect 29472 14940 29500 14980
rect 30466 14968 30472 14980
rect 30524 14968 30530 15020
rect 31386 14968 31392 15020
rect 31444 15017 31450 15020
rect 31680 15017 31708 15048
rect 31444 14971 31456 15017
rect 31665 15011 31723 15017
rect 31665 14977 31677 15011
rect 31711 14977 31723 15011
rect 31665 14971 31723 14977
rect 31444 14968 31450 14971
rect 29012 14912 29500 14940
rect 29546 14900 29552 14952
rect 29604 14940 29610 14952
rect 29733 14943 29791 14949
rect 29733 14940 29745 14943
rect 29604 14912 29745 14940
rect 29604 14900 29610 14912
rect 29733 14909 29745 14912
rect 29779 14909 29791 14943
rect 29733 14903 29791 14909
rect 28920 14872 28948 14900
rect 30285 14875 30343 14881
rect 30285 14872 30297 14875
rect 28920 14844 30297 14872
rect 30285 14841 30297 14844
rect 30331 14841 30343 14875
rect 30285 14835 30343 14841
rect 23845 14807 23903 14813
rect 23845 14804 23857 14807
rect 23768 14776 23857 14804
rect 23661 14767 23719 14773
rect 23845 14773 23857 14776
rect 23891 14773 23903 14807
rect 23845 14767 23903 14773
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 25314 14804 25320 14816
rect 23992 14776 25320 14804
rect 23992 14764 23998 14776
rect 25314 14764 25320 14776
rect 25372 14764 25378 14816
rect 25501 14807 25559 14813
rect 25501 14773 25513 14807
rect 25547 14804 25559 14807
rect 25682 14804 25688 14816
rect 25547 14776 25688 14804
rect 25547 14773 25559 14776
rect 25501 14767 25559 14773
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 26602 14764 26608 14816
rect 26660 14804 26666 14816
rect 27341 14807 27399 14813
rect 27341 14804 27353 14807
rect 26660 14776 27353 14804
rect 26660 14764 26666 14776
rect 27341 14773 27353 14776
rect 27387 14804 27399 14807
rect 27522 14804 27528 14816
rect 27387 14776 27528 14804
rect 27387 14773 27399 14776
rect 27341 14767 27399 14773
rect 27522 14764 27528 14776
rect 27580 14764 27586 14816
rect 28166 14764 28172 14816
rect 28224 14764 28230 14816
rect 29638 14764 29644 14816
rect 29696 14764 29702 14816
rect 29822 14764 29828 14816
rect 29880 14764 29886 14816
rect 1104 14714 32476 14736
rect 1104 14662 4871 14714
rect 4923 14662 4935 14714
rect 4987 14662 4999 14714
rect 5051 14662 5063 14714
rect 5115 14662 5127 14714
rect 5179 14662 12713 14714
rect 12765 14662 12777 14714
rect 12829 14662 12841 14714
rect 12893 14662 12905 14714
rect 12957 14662 12969 14714
rect 13021 14662 20555 14714
rect 20607 14662 20619 14714
rect 20671 14662 20683 14714
rect 20735 14662 20747 14714
rect 20799 14662 20811 14714
rect 20863 14662 28397 14714
rect 28449 14662 28461 14714
rect 28513 14662 28525 14714
rect 28577 14662 28589 14714
rect 28641 14662 28653 14714
rect 28705 14662 32476 14714
rect 1104 14640 32476 14662
rect 3142 14600 3148 14612
rect 2700 14572 3148 14600
rect 2700 14473 2728 14572
rect 3142 14560 3148 14572
rect 3200 14600 3206 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3200 14572 4169 14600
rect 3200 14560 3206 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 8294 14560 8300 14612
rect 8352 14560 8358 14612
rect 8386 14560 8392 14612
rect 8444 14560 8450 14612
rect 9950 14560 9956 14612
rect 10008 14560 10014 14612
rect 10505 14603 10563 14609
rect 10505 14569 10517 14603
rect 10551 14600 10563 14603
rect 10778 14600 10784 14612
rect 10551 14572 10784 14600
rect 10551 14569 10563 14572
rect 10505 14563 10563 14569
rect 6362 14492 6368 14544
rect 6420 14532 6426 14544
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 6420 14504 6469 14532
rect 6420 14492 6426 14504
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 8312 14532 8340 14560
rect 8312 14504 8616 14532
rect 6457 14495 6515 14501
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14433 2743 14467
rect 2685 14427 2743 14433
rect 7650 14424 7656 14476
rect 7708 14424 7714 14476
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 8294 14464 8300 14476
rect 7883 14436 8300 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8588 14464 8616 14504
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 10520 14532 10548 14563
rect 10778 14560 10784 14572
rect 10836 14600 10842 14612
rect 12066 14600 12072 14612
rect 10836 14572 12072 14600
rect 10836 14560 10842 14572
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 12710 14560 12716 14612
rect 12768 14560 12774 14612
rect 13265 14603 13323 14609
rect 13265 14569 13277 14603
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 9824 14504 10548 14532
rect 9824 14492 9830 14504
rect 8588 14436 9904 14464
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2593 14399 2651 14405
rect 2593 14396 2605 14399
rect 2464 14368 2605 14396
rect 2464 14356 2470 14368
rect 2593 14365 2605 14368
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 7098 14396 7104 14408
rect 6779 14368 7104 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7668 14396 7696 14424
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7668 14368 7757 14396
rect 7745 14365 7757 14368
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8588 14405 8616 14436
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8168 14368 8401 14396
rect 8168 14356 8174 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14396 9551 14399
rect 9582 14396 9588 14408
rect 9539 14368 9588 14396
rect 9539 14365 9551 14368
rect 9493 14359 9551 14365
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 3973 14331 4031 14337
rect 3973 14328 3985 14331
rect 3568 14300 3985 14328
rect 3568 14288 3574 14300
rect 3973 14297 3985 14300
rect 4019 14297 4031 14331
rect 3973 14291 4031 14297
rect 6457 14331 6515 14337
rect 6457 14297 6469 14331
rect 6503 14328 6515 14331
rect 7650 14328 7656 14340
rect 6503 14300 7656 14328
rect 6503 14297 6515 14300
rect 6457 14291 6515 14297
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 9508 14328 9536 14359
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 9766 14356 9772 14408
rect 9824 14356 9830 14408
rect 9876 14396 9904 14436
rect 11882 14424 11888 14476
rect 11940 14424 11946 14476
rect 13280 14464 13308 14563
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 13504 14572 13553 14600
rect 13504 14560 13510 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 14642 14600 14648 14612
rect 13541 14563 13599 14569
rect 14292 14572 14648 14600
rect 14182 14464 14188 14476
rect 13280 14436 14188 14464
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14292 14473 14320 14572
rect 14642 14560 14648 14572
rect 14700 14600 14706 14612
rect 21177 14603 21235 14609
rect 21177 14600 21189 14603
rect 14700 14572 16896 14600
rect 14700 14560 14706 14572
rect 16868 14473 16896 14572
rect 18616 14572 21189 14600
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14433 14335 14467
rect 14277 14427 14335 14433
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 12437 14399 12495 14405
rect 9876 14368 11560 14396
rect 11422 14328 11428 14340
rect 9508 14300 11428 14328
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 2961 14263 3019 14269
rect 2961 14229 2973 14263
rect 3007 14260 3019 14263
rect 3050 14260 3056 14272
rect 3007 14232 3056 14260
rect 3007 14229 3019 14232
rect 2961 14223 3019 14229
rect 3050 14220 3056 14232
rect 3108 14260 3114 14272
rect 3418 14260 3424 14272
rect 3108 14232 3424 14260
rect 3108 14220 3114 14232
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 4173 14263 4231 14269
rect 4173 14260 4185 14263
rect 3752 14232 4185 14260
rect 3752 14220 3758 14232
rect 4173 14229 4185 14232
rect 4219 14229 4231 14263
rect 4173 14223 4231 14229
rect 4341 14263 4399 14269
rect 4341 14229 4353 14263
rect 4387 14260 4399 14263
rect 4430 14260 4436 14272
rect 4387 14232 4436 14260
rect 4387 14229 4399 14232
rect 4341 14223 4399 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7377 14263 7435 14269
rect 7377 14260 7389 14263
rect 6788 14232 7389 14260
rect 6788 14220 6794 14232
rect 7377 14229 7389 14232
rect 7423 14229 7435 14263
rect 7377 14223 7435 14229
rect 9585 14263 9643 14269
rect 9585 14229 9597 14263
rect 9631 14260 9643 14263
rect 9674 14260 9680 14272
rect 9631 14232 9680 14260
rect 9631 14229 9643 14232
rect 9585 14223 9643 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 11532 14260 11560 14368
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 12483 14368 13124 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 11606 14288 11612 14340
rect 11664 14337 11670 14340
rect 11664 14291 11676 14337
rect 11664 14288 11670 14291
rect 12710 14288 12716 14340
rect 12768 14288 12774 14340
rect 13096 14328 13124 14368
rect 13170 14356 13176 14408
rect 13228 14356 13234 14408
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 13403 14368 14136 14396
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 13630 14328 13636 14340
rect 13096 14300 13636 14328
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 14108 14328 14136 14368
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14533 14399 14591 14405
rect 14533 14396 14545 14399
rect 14424 14368 14545 14396
rect 14424 14356 14430 14368
rect 14533 14365 14545 14368
rect 14579 14365 14591 14399
rect 14533 14359 14591 14365
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15436 14368 16129 14396
rect 15436 14356 15442 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 16132 14328 16160 14359
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 17109 14399 17167 14405
rect 17109 14396 17121 14399
rect 16356 14368 17121 14396
rect 16356 14356 16362 14368
rect 17109 14365 17121 14368
rect 17155 14365 17167 14399
rect 17109 14359 17167 14365
rect 18616 14328 18644 14572
rect 21177 14569 21189 14572
rect 21223 14600 21235 14603
rect 21726 14600 21732 14612
rect 21223 14572 21732 14600
rect 21223 14569 21235 14572
rect 21177 14563 21235 14569
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 21818 14560 21824 14612
rect 21876 14600 21882 14612
rect 23290 14600 23296 14612
rect 21876 14572 23296 14600
rect 21876 14560 21882 14572
rect 23290 14560 23296 14572
rect 23348 14560 23354 14612
rect 24302 14560 24308 14612
rect 24360 14600 24366 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24360 14572 24777 14600
rect 24360 14560 24366 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 24765 14563 24823 14569
rect 25130 14560 25136 14612
rect 25188 14560 25194 14612
rect 25222 14560 25228 14612
rect 25280 14600 25286 14612
rect 26234 14600 26240 14612
rect 25280 14572 26240 14600
rect 25280 14560 25286 14572
rect 22186 14424 22192 14476
rect 22244 14464 22250 14476
rect 22554 14464 22560 14476
rect 22244 14436 22560 14464
rect 22244 14424 22250 14436
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 23106 14424 23112 14476
rect 23164 14464 23170 14476
rect 25774 14464 25780 14476
rect 23164 14436 25780 14464
rect 23164 14424 23170 14436
rect 19794 14356 19800 14408
rect 19852 14356 19858 14408
rect 20064 14399 20122 14405
rect 20064 14365 20076 14399
rect 20110 14396 20122 14399
rect 20346 14396 20352 14408
rect 20110 14368 20352 14396
rect 20110 14365 20122 14368
rect 20064 14359 20122 14365
rect 20346 14356 20352 14368
rect 20404 14356 20410 14408
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 22646 14356 22652 14408
rect 22704 14356 22710 14408
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23661 14399 23719 14405
rect 23247 14368 23612 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 14108 14300 15976 14328
rect 16132 14300 18644 14328
rect 15948 14272 15976 14300
rect 18782 14288 18788 14340
rect 18840 14328 18846 14340
rect 23216 14328 23244 14359
rect 18840 14300 23244 14328
rect 18840 14288 18846 14300
rect 12434 14260 12440 14272
rect 11532 14232 12440 14260
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 12529 14263 12587 14269
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 13814 14260 13820 14272
rect 12575 14232 13820 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 15657 14263 15715 14269
rect 15657 14260 15669 14263
rect 15344 14232 15669 14260
rect 15344 14220 15350 14232
rect 15657 14229 15669 14232
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 15988 14232 16313 14260
rect 15988 14220 15994 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 18230 14260 18236 14272
rect 17460 14232 18236 14260
rect 17460 14220 17466 14232
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18966 14220 18972 14272
rect 19024 14260 19030 14272
rect 21818 14260 21824 14272
rect 19024 14232 21824 14260
rect 19024 14220 19030 14232
rect 21818 14220 21824 14232
rect 21876 14220 21882 14272
rect 23584 14260 23612 14368
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 23676 14328 23704 14359
rect 24394 14356 24400 14408
rect 24452 14396 24458 14408
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 24452 14368 24777 14396
rect 24452 14356 24458 14368
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 24946 14356 24952 14408
rect 25004 14356 25010 14408
rect 25130 14356 25136 14408
rect 25188 14396 25194 14408
rect 25701 14405 25729 14436
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 25593 14399 25651 14405
rect 25593 14396 25605 14399
rect 25188 14368 25605 14396
rect 25188 14356 25194 14368
rect 25593 14365 25605 14368
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25686 14399 25744 14405
rect 25686 14365 25698 14399
rect 25732 14365 25744 14399
rect 25686 14359 25744 14365
rect 25866 14356 25872 14408
rect 25924 14356 25930 14408
rect 26077 14399 26135 14405
rect 26077 14365 26089 14399
rect 26123 14396 26135 14399
rect 26165 14396 26193 14572
rect 26234 14560 26240 14572
rect 26292 14560 26298 14612
rect 26881 14603 26939 14609
rect 26881 14569 26893 14603
rect 26927 14600 26939 14603
rect 28166 14600 28172 14612
rect 26927 14572 28172 14600
rect 26927 14569 26939 14572
rect 26881 14563 26939 14569
rect 28166 14560 28172 14572
rect 28224 14560 28230 14612
rect 31110 14600 31116 14612
rect 29748 14572 31116 14600
rect 26326 14492 26332 14544
rect 26384 14532 26390 14544
rect 26384 14504 27016 14532
rect 26384 14492 26390 14504
rect 26602 14424 26608 14476
rect 26660 14464 26666 14476
rect 26988 14473 27016 14504
rect 26789 14467 26847 14473
rect 26789 14464 26801 14467
rect 26660 14436 26801 14464
rect 26660 14424 26666 14436
rect 26789 14433 26801 14436
rect 26835 14433 26847 14467
rect 26789 14427 26847 14433
rect 26973 14467 27031 14473
rect 26973 14433 26985 14467
rect 27019 14433 27031 14467
rect 26973 14427 27031 14433
rect 27706 14424 27712 14476
rect 27764 14464 27770 14476
rect 28810 14464 28816 14476
rect 27764 14436 28816 14464
rect 27764 14424 27770 14436
rect 28810 14424 28816 14436
rect 28868 14464 28874 14476
rect 29748 14473 29776 14572
rect 31110 14560 31116 14572
rect 31168 14560 31174 14612
rect 29733 14467 29791 14473
rect 29733 14464 29745 14467
rect 28868 14436 29745 14464
rect 28868 14424 28874 14436
rect 29733 14433 29745 14436
rect 29779 14433 29791 14467
rect 29733 14427 29791 14433
rect 26123 14368 26193 14396
rect 26123 14365 26135 14368
rect 26077 14359 26135 14365
rect 26234 14356 26240 14408
rect 26292 14396 26298 14408
rect 26697 14399 26755 14405
rect 26697 14396 26709 14399
rect 26292 14368 26709 14396
rect 26292 14356 26298 14368
rect 26697 14365 26709 14368
rect 26743 14365 26755 14399
rect 26697 14359 26755 14365
rect 27430 14356 27436 14408
rect 27488 14396 27494 14408
rect 28261 14399 28319 14405
rect 28261 14396 28273 14399
rect 27488 14368 28273 14396
rect 27488 14356 27494 14368
rect 28261 14365 28273 14368
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28902 14356 28908 14408
rect 28960 14356 28966 14408
rect 29822 14356 29828 14408
rect 29880 14396 29886 14408
rect 29989 14399 30047 14405
rect 29989 14396 30001 14399
rect 29880 14368 30001 14396
rect 29880 14356 29886 14368
rect 29989 14365 30001 14368
rect 30035 14365 30047 14399
rect 29989 14359 30047 14365
rect 25406 14328 25412 14340
rect 23676 14300 25412 14328
rect 25406 14288 25412 14300
rect 25464 14288 25470 14340
rect 25958 14288 25964 14340
rect 26016 14288 26022 14340
rect 28810 14288 28816 14340
rect 28868 14288 28874 14340
rect 30098 14328 30104 14340
rect 28966 14300 30104 14328
rect 23842 14260 23848 14272
rect 23584 14232 23848 14260
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 24210 14220 24216 14272
rect 24268 14260 24274 14272
rect 24946 14260 24952 14272
rect 24268 14232 24952 14260
rect 24268 14220 24274 14232
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 25314 14220 25320 14272
rect 25372 14260 25378 14272
rect 26142 14260 26148 14272
rect 25372 14232 26148 14260
rect 25372 14220 25378 14232
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 26234 14220 26240 14272
rect 26292 14220 26298 14272
rect 28074 14220 28080 14272
rect 28132 14220 28138 14272
rect 28718 14220 28724 14272
rect 28776 14260 28782 14272
rect 28966 14260 28994 14300
rect 30098 14288 30104 14300
rect 30156 14288 30162 14340
rect 28776 14232 28994 14260
rect 28776 14220 28782 14232
rect 29730 14220 29736 14272
rect 29788 14260 29794 14272
rect 31113 14263 31171 14269
rect 31113 14260 31125 14263
rect 29788 14232 31125 14260
rect 29788 14220 29794 14232
rect 31113 14229 31125 14232
rect 31159 14229 31171 14263
rect 31113 14223 31171 14229
rect 1104 14170 32632 14192
rect 1104 14118 8792 14170
rect 8844 14118 8856 14170
rect 8908 14118 8920 14170
rect 8972 14118 8984 14170
rect 9036 14118 9048 14170
rect 9100 14118 16634 14170
rect 16686 14118 16698 14170
rect 16750 14118 16762 14170
rect 16814 14118 16826 14170
rect 16878 14118 16890 14170
rect 16942 14118 24476 14170
rect 24528 14118 24540 14170
rect 24592 14118 24604 14170
rect 24656 14118 24668 14170
rect 24720 14118 24732 14170
rect 24784 14118 32318 14170
rect 32370 14118 32382 14170
rect 32434 14118 32446 14170
rect 32498 14118 32510 14170
rect 32562 14118 32574 14170
rect 32626 14118 32632 14170
rect 1104 14096 32632 14118
rect 3510 14056 3516 14068
rect 2608 14028 3516 14056
rect 2608 13929 2636 14028
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 10502 14056 10508 14068
rect 9732 14028 10508 14056
rect 9732 14016 9738 14028
rect 10502 14016 10508 14028
rect 10560 14056 10566 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10560 14028 10609 14056
rect 10560 14016 10566 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 10597 14019 10655 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 11701 14059 11759 14065
rect 11701 14056 11713 14059
rect 11664 14028 11713 14056
rect 11664 14016 11670 14028
rect 11701 14025 11713 14028
rect 11747 14025 11759 14059
rect 11701 14019 11759 14025
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 13265 14059 13323 14065
rect 13265 14056 13277 14059
rect 12768 14028 13277 14056
rect 12768 14016 12774 14028
rect 13265 14025 13277 14028
rect 13311 14025 13323 14059
rect 13265 14019 13323 14025
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14826 14056 14832 14068
rect 14139 14028 14832 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 3694 13988 3700 14000
rect 3252 13960 3700 13988
rect 3252 13929 3280 13960
rect 3694 13948 3700 13960
rect 3752 13948 3758 14000
rect 5626 13948 5632 14000
rect 5684 13948 5690 14000
rect 5845 13991 5903 13997
rect 5845 13957 5857 13991
rect 5891 13988 5903 13991
rect 6730 13988 6736 14000
rect 5891 13960 6736 13988
rect 5891 13957 5903 13960
rect 5845 13951 5903 13957
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 7800 13960 8217 13988
rect 7800 13948 7806 13960
rect 8205 13957 8217 13960
rect 8251 13957 8263 13991
rect 8205 13951 8263 13957
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 1995 13892 2605 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 1780 13852 1808 13883
rect 3418 13880 3424 13932
rect 3476 13880 3482 13932
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 3602 13880 3608 13932
rect 3660 13880 3666 13932
rect 4522 13880 4528 13932
rect 4580 13880 4586 13932
rect 5644 13920 5672 13948
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 5644 13892 7021 13920
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 9214 13880 9220 13932
rect 9272 13880 9278 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9473 13923 9531 13929
rect 9473 13920 9485 13923
rect 9364 13892 9485 13920
rect 9364 13880 9370 13892
rect 9473 13889 9485 13892
rect 9519 13889 9531 13923
rect 9473 13883 9531 13889
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 11885 13923 11943 13929
rect 11885 13920 11897 13923
rect 10744 13892 11897 13920
rect 10744 13880 10750 13892
rect 11885 13889 11897 13892
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13814 13920 13820 13932
rect 13587 13892 13820 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13814 13880 13820 13892
rect 13872 13920 13878 13932
rect 14108 13920 14136 14019
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 16209 14059 16267 14065
rect 16209 14056 16221 14059
rect 15620 14028 16221 14056
rect 15620 14016 15626 14028
rect 16209 14025 16221 14028
rect 16255 14025 16267 14059
rect 16209 14019 16267 14025
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 23382 14056 23388 14068
rect 18472 14028 23388 14056
rect 18472 14016 18478 14028
rect 23382 14016 23388 14028
rect 23440 14056 23446 14068
rect 26050 14056 26056 14068
rect 23440 14028 26056 14056
rect 23440 14016 23446 14028
rect 26050 14016 26056 14028
rect 26108 14016 26114 14068
rect 31754 14056 31760 14068
rect 26896 14028 31760 14056
rect 15286 13988 15292 14000
rect 14292 13960 15292 13988
rect 14292 13929 14320 13960
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 15841 13991 15899 13997
rect 15841 13957 15853 13991
rect 15887 13988 15899 13991
rect 16114 13988 16120 14000
rect 15887 13960 16120 13988
rect 15887 13957 15899 13960
rect 15841 13951 15899 13957
rect 16114 13948 16120 13960
rect 16172 13948 16178 14000
rect 19705 13991 19763 13997
rect 19705 13957 19717 13991
rect 19751 13988 19763 13991
rect 26896 13988 26924 14028
rect 31754 14016 31760 14028
rect 31812 14016 31818 14068
rect 19751 13960 26924 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 28902 13948 28908 14000
rect 28960 13988 28966 14000
rect 30285 13991 30343 13997
rect 30285 13988 30297 13991
rect 28960 13960 30297 13988
rect 28960 13948 28966 13960
rect 30285 13957 30297 13960
rect 30331 13957 30343 13991
rect 30285 13951 30343 13957
rect 30466 13948 30472 14000
rect 30524 13997 30530 14000
rect 30524 13991 30543 13997
rect 30531 13957 30543 13991
rect 30524 13951 30543 13957
rect 30524 13948 30530 13951
rect 13872 13892 14136 13920
rect 14277 13923 14335 13929
rect 13872 13880 13878 13892
rect 14277 13889 14289 13923
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15378 13920 15384 13932
rect 15059 13892 15384 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 15712 13892 15761 13920
rect 15712 13880 15718 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 17034 13920 17040 13932
rect 16071 13892 17040 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17310 13880 17316 13932
rect 17368 13880 17374 13932
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21784 13892 22017 13920
rect 21784 13880 21790 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 22244 13892 22477 13920
rect 22244 13880 22250 13892
rect 22465 13889 22477 13892
rect 22511 13889 22523 13923
rect 23106 13920 23112 13932
rect 22465 13883 22523 13889
rect 22848 13892 23112 13920
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 1780 13824 2789 13852
rect 2777 13821 2789 13824
rect 2823 13852 2835 13855
rect 3620 13852 3648 13880
rect 2823 13824 3648 13852
rect 3881 13855 3939 13861
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 4246 13852 4252 13864
rect 3927 13824 4252 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4430 13812 4436 13864
rect 4488 13812 4494 13864
rect 4540 13852 4568 13880
rect 13265 13855 13323 13861
rect 4540 13824 5856 13852
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2222 13716 2228 13728
rect 1995 13688 2228 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 2406 13676 2412 13728
rect 2464 13676 2470 13728
rect 4801 13719 4859 13725
rect 4801 13685 4813 13719
rect 4847 13716 4859 13719
rect 5350 13716 5356 13728
rect 4847 13688 5356 13716
rect 4847 13685 4859 13688
rect 4801 13679 4859 13685
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 5828 13725 5856 13824
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13354 13852 13360 13864
rect 13311 13824 13360 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 13449 13855 13507 13861
rect 13449 13821 13461 13855
rect 13495 13852 13507 13855
rect 13630 13852 13636 13864
rect 13495 13824 13636 13852
rect 13495 13821 13507 13824
rect 13449 13815 13507 13821
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15286 13852 15292 13864
rect 15151 13824 15292 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 20438 13852 20444 13864
rect 18288 13824 20444 13852
rect 18288 13812 18294 13824
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 21910 13812 21916 13864
rect 21968 13852 21974 13864
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 21968 13824 22293 13852
rect 21968 13812 21974 13824
rect 22281 13821 22293 13824
rect 22327 13821 22339 13855
rect 22281 13815 22339 13821
rect 22370 13812 22376 13864
rect 22428 13852 22434 13864
rect 22848 13852 22876 13892
rect 23106 13880 23112 13892
rect 23164 13920 23170 13932
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 23164 13892 23213 13920
rect 23164 13880 23170 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23293 13923 23351 13929
rect 23293 13889 23305 13923
rect 23339 13889 23351 13923
rect 23293 13883 23351 13889
rect 22428 13824 22876 13852
rect 22428 13812 22434 13824
rect 22922 13812 22928 13864
rect 22980 13852 22986 13864
rect 23308 13852 23336 13883
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 24489 13923 24547 13929
rect 24489 13920 24501 13923
rect 24452 13892 24501 13920
rect 24452 13880 24458 13892
rect 24489 13889 24501 13892
rect 24535 13889 24547 13923
rect 24489 13883 24547 13889
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25406 13880 25412 13932
rect 25464 13920 25470 13932
rect 25685 13923 25743 13929
rect 25685 13920 25697 13923
rect 25464 13892 25697 13920
rect 25464 13880 25470 13892
rect 25685 13889 25697 13892
rect 25731 13920 25743 13923
rect 26421 13923 26479 13929
rect 26421 13920 26433 13923
rect 25731 13892 26433 13920
rect 25731 13889 25743 13892
rect 25685 13883 25743 13889
rect 26421 13889 26433 13892
rect 26467 13889 26479 13923
rect 26421 13883 26479 13889
rect 26510 13880 26516 13932
rect 26568 13880 26574 13932
rect 27706 13880 27712 13932
rect 27764 13880 27770 13932
rect 27798 13880 27804 13932
rect 27856 13920 27862 13932
rect 27965 13923 28023 13929
rect 27965 13920 27977 13923
rect 27856 13892 27977 13920
rect 27856 13880 27862 13892
rect 27965 13889 27977 13892
rect 28011 13889 28023 13923
rect 27965 13883 28023 13889
rect 29362 13880 29368 13932
rect 29420 13920 29426 13932
rect 29549 13923 29607 13929
rect 29549 13920 29561 13923
rect 29420 13892 29561 13920
rect 29420 13880 29426 13892
rect 29549 13889 29561 13892
rect 29595 13889 29607 13923
rect 29549 13883 29607 13889
rect 29730 13880 29736 13932
rect 29788 13880 29794 13932
rect 29825 13923 29883 13929
rect 29825 13889 29837 13923
rect 29871 13920 29883 13923
rect 30484 13920 30512 13948
rect 31113 13923 31171 13929
rect 31113 13920 31125 13923
rect 29871 13892 30512 13920
rect 30668 13892 31125 13920
rect 29871 13889 29883 13892
rect 29825 13883 29883 13889
rect 22980 13824 23336 13852
rect 22980 13812 22986 13824
rect 24302 13812 24308 13864
rect 24360 13852 24366 13864
rect 24360 13824 24440 13852
rect 24360 13812 24366 13824
rect 6730 13744 6736 13796
rect 6788 13744 6794 13796
rect 17770 13784 17776 13796
rect 14752 13756 17776 13784
rect 14752 13728 14780 13756
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 22940 13784 22968 13812
rect 24412 13793 24440 13824
rect 25038 13812 25044 13864
rect 25096 13852 25102 13864
rect 25501 13855 25559 13861
rect 25501 13852 25513 13855
rect 25096 13824 25513 13852
rect 25096 13812 25102 13824
rect 25501 13821 25513 13824
rect 25547 13821 25559 13855
rect 25501 13815 25559 13821
rect 25866 13812 25872 13864
rect 25924 13852 25930 13864
rect 26694 13852 26700 13864
rect 25924 13824 26700 13852
rect 25924 13812 25930 13824
rect 26694 13812 26700 13824
rect 26752 13812 26758 13864
rect 29638 13852 29644 13864
rect 29564 13824 29644 13852
rect 22480 13756 22968 13784
rect 24397 13787 24455 13793
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13685 5871 13719
rect 5813 13679 5871 13685
rect 5994 13676 6000 13728
rect 6052 13676 6058 13728
rect 6546 13676 6552 13728
rect 6604 13676 6610 13728
rect 8110 13676 8116 13728
rect 8168 13676 8174 13728
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 14734 13716 14740 13728
rect 12676 13688 14740 13716
rect 12676 13676 12682 13688
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 14829 13719 14887 13725
rect 14829 13685 14841 13719
rect 14875 13716 14887 13719
rect 14918 13716 14924 13728
rect 14875 13688 14924 13716
rect 14875 13685 14887 13688
rect 14829 13679 14887 13685
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 15838 13716 15844 13728
rect 15344 13688 15844 13716
rect 15344 13676 15350 13688
rect 15838 13676 15844 13688
rect 15896 13716 15902 13728
rect 17402 13716 17408 13728
rect 15896 13688 17408 13716
rect 15896 13676 15902 13688
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17494 13676 17500 13728
rect 17552 13676 17558 13728
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 22480 13725 22508 13756
rect 24397 13753 24409 13787
rect 24443 13753 24455 13787
rect 26602 13784 26608 13796
rect 24397 13747 24455 13753
rect 25240 13756 26608 13784
rect 22465 13719 22523 13725
rect 22465 13716 22477 13719
rect 22428 13688 22477 13716
rect 22428 13676 22434 13688
rect 22465 13685 22477 13688
rect 22511 13685 22523 13719
rect 22465 13679 22523 13685
rect 22646 13676 22652 13728
rect 22704 13676 22710 13728
rect 24210 13676 24216 13728
rect 24268 13716 24274 13728
rect 24305 13719 24363 13725
rect 24305 13716 24317 13719
rect 24268 13688 24317 13716
rect 24268 13676 24274 13688
rect 24305 13685 24317 13688
rect 24351 13716 24363 13719
rect 25240 13716 25268 13756
rect 26602 13744 26608 13756
rect 26660 13744 26666 13796
rect 29564 13793 29592 13824
rect 29638 13812 29644 13824
rect 29696 13812 29702 13864
rect 30668 13793 30696 13892
rect 31113 13889 31125 13892
rect 31159 13889 31171 13923
rect 31113 13883 31171 13889
rect 31386 13852 31392 13864
rect 31312 13824 31392 13852
rect 31312 13793 31340 13824
rect 31386 13812 31392 13824
rect 31444 13812 31450 13864
rect 29549 13787 29607 13793
rect 29549 13753 29561 13787
rect 29595 13753 29607 13787
rect 29549 13747 29607 13753
rect 30653 13787 30711 13793
rect 30653 13753 30665 13787
rect 30699 13753 30711 13787
rect 30653 13747 30711 13753
rect 31297 13787 31355 13793
rect 31297 13753 31309 13787
rect 31343 13753 31355 13787
rect 31297 13747 31355 13753
rect 24351 13688 25268 13716
rect 24351 13685 24363 13688
rect 24305 13679 24363 13685
rect 25314 13676 25320 13728
rect 25372 13676 25378 13728
rect 25866 13676 25872 13728
rect 25924 13676 25930 13728
rect 29086 13676 29092 13728
rect 29144 13676 29150 13728
rect 30374 13676 30380 13728
rect 30432 13716 30438 13728
rect 30469 13719 30527 13725
rect 30469 13716 30481 13719
rect 30432 13688 30481 13716
rect 30432 13676 30438 13688
rect 30469 13685 30481 13688
rect 30515 13685 30527 13719
rect 30469 13679 30527 13685
rect 1104 13626 32476 13648
rect 1104 13574 4871 13626
rect 4923 13574 4935 13626
rect 4987 13574 4999 13626
rect 5051 13574 5063 13626
rect 5115 13574 5127 13626
rect 5179 13574 12713 13626
rect 12765 13574 12777 13626
rect 12829 13574 12841 13626
rect 12893 13574 12905 13626
rect 12957 13574 12969 13626
rect 13021 13574 20555 13626
rect 20607 13574 20619 13626
rect 20671 13574 20683 13626
rect 20735 13574 20747 13626
rect 20799 13574 20811 13626
rect 20863 13574 28397 13626
rect 28449 13574 28461 13626
rect 28513 13574 28525 13626
rect 28577 13574 28589 13626
rect 28641 13574 28653 13626
rect 28705 13574 32476 13626
rect 1104 13552 32476 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 3108 13484 4169 13512
rect 3108 13472 3114 13484
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 5353 13515 5411 13521
rect 5353 13481 5365 13515
rect 5399 13512 5411 13515
rect 5902 13512 5908 13524
rect 5399 13484 5908 13512
rect 5399 13481 5411 13484
rect 5353 13475 5411 13481
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 7098 13472 7104 13524
rect 7156 13472 7162 13524
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 8168 13484 9628 13512
rect 8168 13472 8174 13484
rect 3421 13447 3479 13453
rect 3421 13413 3433 13447
rect 3467 13444 3479 13447
rect 4341 13447 4399 13453
rect 3467 13416 4200 13444
rect 3467 13413 3479 13416
rect 3421 13407 3479 13413
rect 2240 13348 4108 13376
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2240 13317 2268 13348
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 2188 13280 2237 13308
rect 2188 13268 2194 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 2682 13268 2688 13320
rect 2740 13268 2746 13320
rect 2884 13317 2912 13348
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 2958 13268 2964 13320
rect 3016 13268 3022 13320
rect 3050 13268 3056 13320
rect 3108 13268 3114 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 3252 13240 3280 13271
rect 2464 13212 3280 13240
rect 2464 13200 2470 13212
rect 3326 13200 3332 13252
rect 3384 13240 3390 13252
rect 3973 13243 4031 13249
rect 3973 13240 3985 13243
rect 3384 13212 3985 13240
rect 3384 13200 3390 13212
rect 3973 13209 3985 13212
rect 4019 13209 4031 13243
rect 4080 13240 4108 13348
rect 4172 13308 4200 13416
rect 4341 13413 4353 13447
rect 4387 13444 4399 13447
rect 9493 13447 9551 13453
rect 4387 13416 6132 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 4304 13348 5181 13376
rect 4304 13336 4310 13348
rect 5169 13345 5181 13348
rect 5215 13345 5227 13379
rect 5169 13339 5227 13345
rect 5994 13336 6000 13388
rect 6052 13336 6058 13388
rect 6104 13385 6132 13416
rect 9493 13413 9505 13447
rect 9539 13413 9551 13447
rect 9600 13444 9628 13484
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 10192 13484 10425 13512
rect 10192 13472 10198 13484
rect 10413 13481 10425 13484
rect 10459 13481 10471 13515
rect 10413 13475 10471 13481
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 10597 13515 10655 13521
rect 10597 13512 10609 13515
rect 10560 13484 10609 13512
rect 10560 13472 10566 13484
rect 10597 13481 10609 13484
rect 10643 13481 10655 13515
rect 12618 13512 12624 13524
rect 10597 13475 10655 13481
rect 10704 13484 12624 13512
rect 10704 13444 10732 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 14642 13512 14648 13524
rect 13004 13484 14648 13512
rect 12897 13447 12955 13453
rect 12897 13444 12909 13447
rect 9600 13416 10732 13444
rect 11256 13416 12909 13444
rect 9493 13407 9551 13413
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13345 6147 13379
rect 9508 13376 9536 13407
rect 6089 13339 6147 13345
rect 6656 13348 9536 13376
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4172 13280 4905 13308
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5350 13268 5356 13320
rect 5408 13268 5414 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 4173 13243 4231 13249
rect 4173 13240 4185 13243
rect 4080 13212 4185 13240
rect 3973 13203 4031 13209
rect 4173 13209 4185 13212
rect 4219 13209 4231 13243
rect 6380 13240 6408 13271
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 6656 13240 6684 13348
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7285 13311 7343 13317
rect 7285 13308 7297 13311
rect 6788 13280 7297 13308
rect 6788 13268 6794 13280
rect 7285 13277 7297 13280
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7558 13268 7564 13320
rect 7616 13268 7622 13320
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 9674 13308 9680 13320
rect 9539 13280 9680 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 4173 13203 4231 13209
rect 4264 13212 6408 13240
rect 6564 13212 6684 13240
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 3234 13172 3240 13184
rect 2179 13144 3240 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4264 13172 4292 13212
rect 3476 13144 4292 13172
rect 3476 13132 3482 13144
rect 5534 13132 5540 13184
rect 5592 13132 5598 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 6273 13175 6331 13181
rect 6273 13172 6285 13175
rect 5868 13144 6285 13172
rect 5868 13132 5874 13144
rect 6273 13141 6285 13144
rect 6319 13172 6331 13175
rect 6564 13172 6592 13212
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7668 13240 7696 13271
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 9766 13268 9772 13320
rect 9824 13268 9830 13320
rect 11256 13317 11284 13416
rect 12897 13413 12909 13416
rect 12943 13413 12955 13447
rect 12897 13407 12955 13413
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 10704 13280 11253 13308
rect 6880 13212 7696 13240
rect 6880 13200 6886 13212
rect 9398 13200 9404 13252
rect 9456 13240 9462 13252
rect 10565 13243 10623 13249
rect 10565 13240 10577 13243
rect 9456 13212 10577 13240
rect 9456 13200 9462 13212
rect 10565 13209 10577 13212
rect 10611 13240 10623 13243
rect 10704 13240 10732 13280
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12158 13268 12164 13320
rect 12216 13268 12222 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13004 13308 13032 13484
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 18785 13515 18843 13521
rect 18785 13512 18797 13515
rect 15436 13484 18797 13512
rect 15436 13472 15442 13484
rect 18785 13481 18797 13484
rect 18831 13512 18843 13515
rect 18966 13512 18972 13524
rect 18831 13484 18972 13512
rect 18831 13481 18843 13484
rect 18785 13475 18843 13481
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 21542 13472 21548 13524
rect 21600 13512 21606 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 21600 13484 22109 13512
rect 21600 13472 21606 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 22204 13484 25728 13512
rect 14090 13444 14096 13456
rect 13096 13416 14096 13444
rect 13096 13317 13124 13416
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 15010 13444 15016 13456
rect 14476 13416 15016 13444
rect 12943 13280 13032 13308
rect 13081 13311 13139 13317
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 14476 13317 14504 13416
rect 15010 13404 15016 13416
rect 15068 13404 15074 13456
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 15470 13444 15476 13456
rect 15252 13416 15476 13444
rect 15252 13404 15258 13416
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 19426 13404 19432 13456
rect 19484 13404 19490 13456
rect 19518 13404 19524 13456
rect 19576 13444 19582 13456
rect 21913 13447 21971 13453
rect 21913 13444 21925 13447
rect 19576 13416 21925 13444
rect 19576 13404 19582 13416
rect 21913 13413 21925 13416
rect 21959 13413 21971 13447
rect 21913 13407 21971 13413
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 10611 13212 10732 13240
rect 10611 13209 10623 13212
rect 10565 13203 10623 13209
rect 10778 13200 10784 13252
rect 10836 13200 10842 13252
rect 14660 13240 14688 13339
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 20165 13379 20223 13385
rect 20165 13376 20177 13379
rect 18472 13348 20177 13376
rect 18472 13336 18478 13348
rect 20165 13345 20177 13348
rect 20211 13345 20223 13379
rect 22204 13376 22232 13484
rect 25593 13447 25651 13453
rect 25593 13444 25605 13447
rect 22756 13416 25605 13444
rect 20165 13339 20223 13345
rect 20272 13348 22232 13376
rect 22281 13379 22339 13385
rect 14734 13268 14740 13320
rect 14792 13268 14798 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 14976 13280 15301 13308
rect 14976 13268 14982 13280
rect 15289 13277 15301 13280
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 15562 13268 15568 13320
rect 15620 13308 15626 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 15620 13280 17417 13308
rect 15620 13268 15626 13280
rect 17405 13277 17417 13280
rect 17451 13277 17463 13311
rect 17405 13271 17463 13277
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17661 13311 17719 13317
rect 17661 13308 17673 13311
rect 17552 13280 17673 13308
rect 17552 13268 17558 13280
rect 17661 13277 17673 13280
rect 17707 13277 17719 13311
rect 17661 13271 17719 13277
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 19751 13280 20208 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 16114 13240 16120 13252
rect 14660 13212 16120 13240
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 17770 13200 17776 13252
rect 17828 13240 17834 13252
rect 20180 13249 20208 13280
rect 19429 13243 19487 13249
rect 19429 13240 19441 13243
rect 17828 13212 19441 13240
rect 17828 13200 17834 13212
rect 19429 13209 19441 13212
rect 19475 13240 19487 13243
rect 20165 13243 20223 13249
rect 19475 13212 20116 13240
rect 19475 13209 19487 13212
rect 19429 13203 19487 13209
rect 6319 13144 6592 13172
rect 6319 13141 6331 13144
rect 6273 13135 6331 13141
rect 6638 13132 6644 13184
rect 6696 13132 6702 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 9364 13144 9689 13172
rect 9364 13132 9370 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 11422 13132 11428 13184
rect 11480 13132 11486 13184
rect 12066 13132 12072 13184
rect 12124 13132 12130 13184
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13504 13144 13553 13172
rect 13504 13132 13510 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 13688 13144 14289 13172
rect 13688 13132 13694 13144
rect 14277 13141 14289 13144
rect 14323 13141 14335 13175
rect 14277 13135 14335 13141
rect 14366 13132 14372 13184
rect 14424 13172 14430 13184
rect 15102 13172 15108 13184
rect 14424 13144 15108 13172
rect 14424 13132 14430 13144
rect 15102 13132 15108 13144
rect 15160 13172 15166 13184
rect 15381 13175 15439 13181
rect 15381 13172 15393 13175
rect 15160 13144 15393 13172
rect 15160 13132 15166 13144
rect 15381 13141 15393 13144
rect 15427 13141 15439 13175
rect 15381 13135 15439 13141
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19576 13144 19625 13172
rect 19576 13132 19582 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 20088 13172 20116 13212
rect 20165 13209 20177 13243
rect 20211 13209 20223 13243
rect 20165 13203 20223 13209
rect 20272 13172 20300 13348
rect 22281 13345 22293 13379
rect 22327 13376 22339 13379
rect 22554 13376 22560 13388
rect 22327 13348 22560 13376
rect 22327 13345 22339 13348
rect 22281 13339 22339 13345
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 20346 13268 20352 13320
rect 20404 13268 20410 13320
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13308 21511 13311
rect 21542 13308 21548 13320
rect 21499 13280 21548 13308
rect 21499 13277 21511 13280
rect 21453 13271 21511 13277
rect 20456 13240 20484 13271
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13308 22155 13311
rect 22756 13308 22784 13416
rect 25593 13413 25605 13416
rect 25639 13413 25651 13447
rect 25700 13444 25728 13484
rect 25958 13472 25964 13524
rect 26016 13472 26022 13524
rect 26326 13512 26332 13524
rect 26068 13484 26332 13512
rect 26068 13444 26096 13484
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 27798 13472 27804 13524
rect 27856 13472 27862 13524
rect 28258 13472 28264 13524
rect 28316 13512 28322 13524
rect 28353 13515 28411 13521
rect 28353 13512 28365 13515
rect 28316 13484 28365 13512
rect 28316 13472 28322 13484
rect 28353 13481 28365 13484
rect 28399 13481 28411 13515
rect 29546 13512 29552 13524
rect 28353 13475 28411 13481
rect 29104 13484 29552 13512
rect 25700 13416 26096 13444
rect 25593 13407 25651 13413
rect 26142 13404 26148 13456
rect 26200 13444 26206 13456
rect 26789 13447 26847 13453
rect 26789 13444 26801 13447
rect 26200 13416 26801 13444
rect 26200 13404 26206 13416
rect 26789 13413 26801 13416
rect 26835 13444 26847 13447
rect 28994 13444 29000 13456
rect 26835 13416 29000 13444
rect 26835 13413 26847 13416
rect 26789 13407 26847 13413
rect 28994 13404 29000 13416
rect 29052 13404 29058 13456
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 24302 13376 24308 13388
rect 23523 13348 24308 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 24302 13336 24308 13348
rect 24360 13336 24366 13388
rect 25961 13379 26019 13385
rect 24780 13348 25912 13376
rect 22143 13280 22784 13308
rect 23385 13311 23443 13317
rect 22143 13277 22155 13280
rect 22097 13271 22155 13277
rect 23385 13277 23397 13311
rect 23431 13277 23443 13311
rect 23385 13271 23443 13277
rect 22112 13240 22140 13271
rect 20456 13212 22140 13240
rect 22557 13243 22615 13249
rect 22557 13209 22569 13243
rect 22603 13209 22615 13243
rect 22557 13203 22615 13209
rect 20088 13144 20300 13172
rect 19613 13135 19671 13141
rect 21358 13132 21364 13184
rect 21416 13132 21422 13184
rect 22572 13172 22600 13203
rect 23290 13200 23296 13252
rect 23348 13240 23354 13252
rect 23400 13240 23428 13271
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 24780 13317 24808 13348
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 24268 13280 24593 13308
rect 24268 13268 24274 13280
rect 24581 13277 24593 13280
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 25314 13268 25320 13320
rect 25372 13308 25378 13320
rect 25777 13311 25835 13317
rect 25777 13308 25789 13311
rect 25372 13280 25789 13308
rect 25372 13268 25378 13280
rect 25777 13277 25789 13280
rect 25823 13277 25835 13311
rect 25884 13308 25912 13348
rect 25961 13345 25973 13379
rect 26007 13376 26019 13379
rect 26234 13376 26240 13388
rect 26007 13348 26240 13376
rect 26007 13345 26019 13348
rect 25961 13339 26019 13345
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 26326 13336 26332 13388
rect 26384 13376 26390 13388
rect 27709 13379 27767 13385
rect 27709 13376 27721 13379
rect 26384 13348 27721 13376
rect 26384 13336 26390 13348
rect 27709 13345 27721 13348
rect 27755 13376 27767 13379
rect 29104 13376 29132 13484
rect 29546 13472 29552 13484
rect 29604 13512 29610 13524
rect 30926 13512 30932 13524
rect 29604 13484 30932 13512
rect 29604 13472 29610 13484
rect 30926 13472 30932 13484
rect 30984 13472 30990 13524
rect 29178 13404 29184 13456
rect 29236 13444 29242 13456
rect 30006 13444 30012 13456
rect 29236 13416 30012 13444
rect 29236 13404 29242 13416
rect 30006 13404 30012 13416
rect 30064 13404 30070 13456
rect 27755 13348 29132 13376
rect 27755 13345 27767 13348
rect 27709 13339 27767 13345
rect 29454 13336 29460 13388
rect 29512 13376 29518 13388
rect 30193 13379 30251 13385
rect 30193 13376 30205 13379
rect 29512 13348 30205 13376
rect 29512 13336 29518 13348
rect 30193 13345 30205 13348
rect 30239 13345 30251 13379
rect 30193 13339 30251 13345
rect 25976 13308 26096 13310
rect 26510 13308 26516 13320
rect 25884 13282 26516 13308
rect 25884 13280 26004 13282
rect 26068 13280 26516 13282
rect 25777 13271 25835 13277
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13308 26755 13311
rect 26786 13308 26792 13320
rect 26743 13280 26792 13308
rect 26743 13277 26755 13280
rect 26697 13271 26755 13277
rect 26786 13268 26792 13280
rect 26844 13268 26850 13320
rect 27614 13268 27620 13320
rect 27672 13268 27678 13320
rect 27798 13268 27804 13320
rect 27856 13308 27862 13320
rect 28261 13311 28319 13317
rect 28261 13308 28273 13311
rect 27856 13280 28273 13308
rect 27856 13268 27862 13280
rect 28261 13277 28273 13280
rect 28307 13277 28319 13311
rect 28261 13271 28319 13277
rect 28445 13311 28503 13317
rect 28445 13277 28457 13311
rect 28491 13308 28503 13311
rect 28718 13308 28724 13320
rect 28491 13280 28724 13308
rect 28491 13277 28503 13280
rect 28445 13271 28503 13277
rect 28718 13268 28724 13280
rect 28776 13268 28782 13320
rect 28905 13311 28963 13317
rect 28905 13277 28917 13311
rect 28951 13308 28963 13311
rect 28994 13308 29000 13320
rect 28951 13280 29000 13308
rect 28951 13277 28963 13280
rect 28905 13271 28963 13277
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 29181 13311 29239 13317
rect 29181 13277 29193 13311
rect 29227 13308 29239 13311
rect 29914 13308 29920 13320
rect 29227 13280 29920 13308
rect 29227 13277 29239 13280
rect 29181 13271 29239 13277
rect 29914 13268 29920 13280
rect 29972 13308 29978 13320
rect 30009 13311 30067 13317
rect 30009 13308 30021 13311
rect 29972 13280 30021 13308
rect 29972 13268 29978 13280
rect 30009 13277 30021 13280
rect 30055 13277 30067 13311
rect 30009 13271 30067 13277
rect 23348 13212 23428 13240
rect 23348 13200 23354 13212
rect 24670 13200 24676 13252
rect 24728 13200 24734 13252
rect 25958 13200 25964 13252
rect 26016 13240 26022 13252
rect 26142 13240 26148 13252
rect 26016 13212 26148 13240
rect 26016 13200 26022 13212
rect 26142 13200 26148 13212
rect 26200 13200 26206 13252
rect 26234 13200 26240 13252
rect 26292 13200 26298 13252
rect 27341 13243 27399 13249
rect 27341 13209 27353 13243
rect 27387 13240 27399 13243
rect 29012 13240 29040 13268
rect 29733 13243 29791 13249
rect 29733 13240 29745 13243
rect 27387 13212 27568 13240
rect 29012 13212 29745 13240
rect 27387 13209 27399 13212
rect 27341 13203 27399 13209
rect 22738 13172 22744 13184
rect 22572 13144 22744 13172
rect 22738 13132 22744 13144
rect 22796 13172 22802 13184
rect 23017 13175 23075 13181
rect 23017 13172 23029 13175
rect 22796 13144 23029 13172
rect 22796 13132 22802 13144
rect 23017 13141 23029 13144
rect 23063 13141 23075 13175
rect 23017 13135 23075 13141
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 27430 13172 27436 13184
rect 23900 13144 27436 13172
rect 23900 13132 23906 13144
rect 27430 13132 27436 13144
rect 27488 13132 27494 13184
rect 27540 13172 27568 13212
rect 29733 13209 29745 13212
rect 29779 13209 29791 13243
rect 29733 13203 29791 13209
rect 27706 13172 27712 13184
rect 27540 13144 27712 13172
rect 27706 13132 27712 13144
rect 27764 13132 27770 13184
rect 27890 13132 27896 13184
rect 27948 13172 27954 13184
rect 28997 13175 29055 13181
rect 28997 13172 29009 13175
rect 27948 13144 29009 13172
rect 27948 13132 27954 13144
rect 28997 13141 29009 13144
rect 29043 13172 29055 13175
rect 29638 13172 29644 13184
rect 29043 13144 29644 13172
rect 29043 13141 29055 13144
rect 28997 13135 29055 13141
rect 29638 13132 29644 13144
rect 29696 13172 29702 13184
rect 29825 13175 29883 13181
rect 29825 13172 29837 13175
rect 29696 13144 29837 13172
rect 29696 13132 29702 13144
rect 29825 13141 29837 13144
rect 29871 13141 29883 13175
rect 29825 13135 29883 13141
rect 1104 13082 32632 13104
rect 1104 13030 8792 13082
rect 8844 13030 8856 13082
rect 8908 13030 8920 13082
rect 8972 13030 8984 13082
rect 9036 13030 9048 13082
rect 9100 13030 16634 13082
rect 16686 13030 16698 13082
rect 16750 13030 16762 13082
rect 16814 13030 16826 13082
rect 16878 13030 16890 13082
rect 16942 13030 24476 13082
rect 24528 13030 24540 13082
rect 24592 13030 24604 13082
rect 24656 13030 24668 13082
rect 24720 13030 24732 13082
rect 24784 13030 32318 13082
rect 32370 13030 32382 13082
rect 32434 13030 32446 13082
rect 32498 13030 32510 13082
rect 32562 13030 32574 13082
rect 32626 13030 32632 13082
rect 1104 13008 32632 13030
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 2869 12971 2927 12977
rect 2869 12968 2881 12971
rect 2740 12940 2881 12968
rect 2740 12928 2746 12940
rect 2869 12937 2881 12940
rect 2915 12937 2927 12971
rect 3970 12968 3976 12980
rect 2869 12931 2927 12937
rect 3160 12940 3976 12968
rect 2317 12903 2375 12909
rect 2317 12869 2329 12903
rect 2363 12900 2375 12903
rect 2363 12872 2774 12900
rect 2363 12869 2375 12872
rect 2317 12863 2375 12869
rect 2222 12792 2228 12844
rect 2280 12792 2286 12844
rect 2406 12792 2412 12844
rect 2464 12792 2470 12844
rect 2746 12764 2774 12872
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 3160 12841 3188 12940
rect 3970 12928 3976 12940
rect 4028 12968 4034 12980
rect 4893 12971 4951 12977
rect 4893 12968 4905 12971
rect 4028 12940 4905 12968
rect 4028 12928 4034 12940
rect 4893 12937 4905 12940
rect 4939 12937 4951 12971
rect 4893 12931 4951 12937
rect 5810 12928 5816 12980
rect 5868 12928 5874 12980
rect 5902 12928 5908 12980
rect 5960 12928 5966 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12937 8171 12971
rect 8113 12931 8171 12937
rect 4062 12860 4068 12912
rect 4120 12909 4126 12912
rect 4120 12903 4183 12909
rect 4120 12869 4137 12903
rect 4171 12869 4183 12903
rect 4120 12863 4183 12869
rect 4341 12903 4399 12909
rect 4341 12869 4353 12903
rect 4387 12900 4399 12903
rect 4430 12900 4436 12912
rect 4387 12872 4436 12900
rect 4387 12869 4399 12872
rect 4341 12863 4399 12869
rect 4120 12860 4126 12863
rect 4430 12860 4436 12872
rect 4488 12900 4494 12912
rect 5721 12903 5779 12909
rect 4488 12872 5028 12900
rect 4488 12860 4494 12872
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 2924 12804 3065 12832
rect 2924 12792 2930 12804
rect 3053 12801 3065 12804
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3234 12792 3240 12844
rect 3292 12792 3298 12844
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3418 12832 3424 12844
rect 3375 12804 3424 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3344 12764 3372 12795
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 3694 12832 3700 12844
rect 3559 12804 3700 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 5000 12841 5028 12872
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 6546 12900 6552 12912
rect 5767 12872 6552 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 8128 12900 8156 12931
rect 9306 12928 9312 12980
rect 9364 12928 9370 12980
rect 15654 12968 15660 12980
rect 15304 12940 15660 12968
rect 12158 12900 12164 12912
rect 6656 12872 12164 12900
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 4985 12835 5043 12841
rect 4847 12804 4916 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 2746 12736 3372 12764
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3142 12696 3148 12708
rect 2924 12668 3148 12696
rect 2924 12656 2930 12668
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 3292 12668 4200 12696
rect 3292 12656 3298 12668
rect 3694 12588 3700 12640
rect 3752 12628 3758 12640
rect 4172 12637 4200 12668
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 3752 12600 3985 12628
rect 3752 12588 3758 12600
rect 3973 12597 3985 12600
rect 4019 12597 4031 12631
rect 3973 12591 4031 12597
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4888 12628 4916 12804
rect 4985 12801 4997 12835
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 5000 12764 5028 12795
rect 5626 12792 5632 12844
rect 5684 12792 5690 12844
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6454 12832 6460 12844
rect 6043 12804 6460 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 6454 12792 6460 12804
rect 6512 12832 6518 12844
rect 6656 12832 6684 12872
rect 12158 12860 12164 12872
rect 12216 12900 12222 12912
rect 14550 12900 14556 12912
rect 12216 12872 14556 12900
rect 12216 12860 12222 12872
rect 14550 12860 14556 12872
rect 14608 12900 14614 12912
rect 15304 12900 15332 12940
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 18322 12928 18328 12980
rect 18380 12928 18386 12980
rect 20346 12928 20352 12980
rect 20404 12968 20410 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 20404 12940 22017 12968
rect 20404 12928 20410 12940
rect 22005 12937 22017 12940
rect 22051 12937 22063 12971
rect 22005 12931 22063 12937
rect 22649 12971 22707 12977
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 23290 12968 23296 12980
rect 22695 12940 23296 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 24670 12968 24676 12980
rect 23716 12940 24676 12968
rect 23716 12928 23722 12940
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25222 12968 25228 12980
rect 25004 12940 25228 12968
rect 25004 12928 25010 12940
rect 25222 12928 25228 12940
rect 25280 12968 25286 12980
rect 25280 12940 26096 12968
rect 25280 12928 25286 12940
rect 14608 12872 15332 12900
rect 14608 12860 14614 12872
rect 7006 12841 7012 12844
rect 6512 12804 6684 12832
rect 6512 12792 6518 12804
rect 7000 12795 7012 12841
rect 7006 12792 7012 12795
rect 7064 12792 7070 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9582 12832 9588 12844
rect 9539 12804 9588 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9858 12832 9864 12844
rect 9723 12804 9864 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 11514 12832 11520 12844
rect 10551 12804 11520 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 13170 12792 13176 12844
rect 13228 12792 13234 12844
rect 13446 12841 13452 12844
rect 13440 12832 13452 12841
rect 13407 12804 13452 12832
rect 13440 12795 13452 12804
rect 13446 12792 13452 12795
rect 13504 12792 13510 12844
rect 13906 12792 13912 12844
rect 13964 12832 13970 12844
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 13964 12804 15025 12832
rect 13964 12792 13970 12804
rect 15013 12801 15025 12804
rect 15059 12801 15071 12835
rect 15013 12795 15071 12801
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15304 12841 15332 12872
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 16114 12900 16120 12912
rect 15427 12872 16120 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 16114 12860 16120 12872
rect 16172 12900 16178 12912
rect 18230 12900 18236 12912
rect 16172 12872 18236 12900
rect 16172 12860 16178 12872
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 19426 12860 19432 12912
rect 19484 12909 19490 12912
rect 19484 12900 19496 12909
rect 19484 12872 19529 12900
rect 19484 12863 19496 12872
rect 19484 12860 19490 12863
rect 20898 12860 20904 12912
rect 20956 12900 20962 12912
rect 20956 12872 23336 12900
rect 20956 12860 20962 12872
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 15160 12804 15209 12832
rect 15160 12792 15166 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15519 12835 15577 12841
rect 15519 12801 15531 12835
rect 15565 12832 15577 12835
rect 16022 12832 16028 12844
rect 15565 12804 16028 12832
rect 15565 12801 15577 12804
rect 15519 12795 15577 12801
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 21192 12841 21220 12872
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12801 21235 12835
rect 21177 12795 21235 12801
rect 21358 12792 21364 12844
rect 21416 12832 21422 12844
rect 22281 12835 22339 12841
rect 22281 12832 22293 12835
rect 21416 12804 22293 12832
rect 21416 12792 21422 12804
rect 22281 12801 22293 12804
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22738 12792 22744 12844
rect 22796 12792 22802 12844
rect 23308 12841 23336 12872
rect 24320 12872 25452 12900
rect 24320 12844 24348 12872
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 23720 12835 23778 12841
rect 23720 12801 23732 12835
rect 23766 12832 23778 12835
rect 23842 12832 23848 12844
rect 23766 12804 23848 12832
rect 23766 12801 23778 12804
rect 23720 12795 23778 12801
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 24302 12792 24308 12844
rect 24360 12792 24366 12844
rect 24489 12835 24547 12841
rect 24489 12801 24501 12835
rect 24535 12801 24547 12835
rect 24489 12795 24547 12801
rect 5718 12764 5724 12776
rect 5000 12736 5724 12764
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 6733 12767 6791 12773
rect 6733 12764 6745 12767
rect 6604 12736 6745 12764
rect 6604 12724 6610 12736
rect 6733 12733 6745 12736
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 10594 12724 10600 12776
rect 10652 12724 10658 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 14568 12736 15669 12764
rect 14458 12656 14464 12708
rect 14516 12696 14522 12708
rect 14568 12705 14596 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 19794 12764 19800 12776
rect 19751 12736 19800 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 19794 12724 19800 12736
rect 19852 12764 19858 12776
rect 20898 12764 20904 12776
rect 19852 12736 20904 12764
rect 19852 12724 19858 12736
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 21453 12767 21511 12773
rect 21453 12733 21465 12767
rect 21499 12764 21511 12767
rect 22094 12764 22100 12776
rect 21499 12736 22100 12764
rect 21499 12733 21511 12736
rect 21453 12727 21511 12733
rect 22094 12724 22100 12736
rect 22152 12724 22158 12776
rect 23198 12724 23204 12776
rect 23256 12724 23262 12776
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 14516 12668 14565 12696
rect 14516 12656 14522 12668
rect 14553 12665 14565 12668
rect 14599 12665 14611 12699
rect 14553 12659 14611 12665
rect 15194 12656 15200 12708
rect 15252 12696 15258 12708
rect 15930 12696 15936 12708
rect 15252 12668 15936 12696
rect 15252 12656 15258 12668
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 21269 12699 21327 12705
rect 21269 12696 21281 12699
rect 20496 12668 21281 12696
rect 20496 12656 20502 12668
rect 21269 12665 21281 12668
rect 21315 12665 21327 12699
rect 21269 12659 21327 12665
rect 21361 12699 21419 12705
rect 21361 12665 21373 12699
rect 21407 12696 21419 12699
rect 22278 12696 22284 12708
rect 21407 12668 22284 12696
rect 21407 12665 21419 12668
rect 21361 12659 21419 12665
rect 7374 12628 7380 12640
rect 4203 12600 7380 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 10226 12588 10232 12640
rect 10284 12588 10290 12640
rect 13538 12588 13544 12640
rect 13596 12628 13602 12640
rect 19518 12628 19524 12640
rect 13596 12600 19524 12628
rect 13596 12588 13602 12600
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 21284 12628 21312 12659
rect 22278 12656 22284 12668
rect 22336 12656 22342 12708
rect 22465 12699 22523 12705
rect 22465 12665 22477 12699
rect 22511 12696 22523 12699
rect 23845 12699 23903 12705
rect 23845 12696 23857 12699
rect 22511 12668 23857 12696
rect 22511 12665 22523 12668
rect 22465 12659 22523 12665
rect 23845 12665 23857 12668
rect 23891 12665 23903 12699
rect 23845 12659 23903 12665
rect 22186 12628 22192 12640
rect 21284 12600 22192 12628
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 22373 12631 22431 12637
rect 22373 12597 22385 12631
rect 22419 12628 22431 12631
rect 22830 12628 22836 12640
rect 22419 12600 22836 12628
rect 22419 12597 22431 12600
rect 22373 12591 22431 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 24504 12628 24532 12795
rect 25424 12696 25452 12872
rect 25498 12860 25504 12912
rect 25556 12900 25562 12912
rect 25961 12903 26019 12909
rect 25961 12900 25973 12903
rect 25556 12872 25973 12900
rect 25556 12860 25562 12872
rect 25961 12869 25973 12872
rect 26007 12869 26019 12903
rect 26068 12900 26096 12940
rect 26142 12928 26148 12980
rect 26200 12968 26206 12980
rect 26329 12971 26387 12977
rect 26329 12968 26341 12971
rect 26200 12940 26341 12968
rect 26200 12928 26206 12940
rect 26329 12937 26341 12940
rect 26375 12937 26387 12971
rect 26329 12931 26387 12937
rect 27430 12928 27436 12980
rect 27488 12968 27494 12980
rect 28994 12968 29000 12980
rect 27488 12940 29000 12968
rect 27488 12928 27494 12940
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 28261 12903 28319 12909
rect 28261 12900 28273 12903
rect 26068 12872 28273 12900
rect 25961 12863 26019 12869
rect 28261 12869 28273 12872
rect 28307 12869 28319 12903
rect 28261 12863 28319 12869
rect 28445 12903 28503 12909
rect 28445 12869 28457 12903
rect 28491 12900 28503 12903
rect 29178 12900 29184 12912
rect 28491 12872 29184 12900
rect 28491 12869 28503 12872
rect 28445 12863 28503 12869
rect 29178 12860 29184 12872
rect 29236 12860 29242 12912
rect 32030 12900 32036 12912
rect 29380 12872 32036 12900
rect 25682 12792 25688 12844
rect 25740 12792 25746 12844
rect 25778 12835 25836 12841
rect 25778 12801 25790 12835
rect 25824 12801 25836 12835
rect 25778 12795 25836 12801
rect 25590 12724 25596 12776
rect 25648 12764 25654 12776
rect 25793 12764 25821 12795
rect 26050 12792 26056 12844
rect 26108 12792 26114 12844
rect 26150 12835 26208 12841
rect 26150 12801 26162 12835
rect 26196 12801 26208 12835
rect 26150 12795 26208 12801
rect 25648 12736 25821 12764
rect 25648 12724 25654 12736
rect 25958 12724 25964 12776
rect 26016 12764 26022 12776
rect 26160 12764 26188 12795
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 27304 12804 27353 12832
rect 27304 12792 27310 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12832 27675 12835
rect 27706 12832 27712 12844
rect 27663 12804 27712 12832
rect 27663 12801 27675 12804
rect 27617 12795 27675 12801
rect 27706 12792 27712 12804
rect 27764 12792 27770 12844
rect 28629 12835 28687 12841
rect 28629 12801 28641 12835
rect 28675 12832 28687 12835
rect 28902 12832 28908 12844
rect 28675 12804 28908 12832
rect 28675 12801 28687 12804
rect 28629 12795 28687 12801
rect 28902 12792 28908 12804
rect 28960 12832 28966 12844
rect 29380 12841 29408 12872
rect 32030 12860 32036 12872
rect 32088 12860 32094 12912
rect 29089 12835 29147 12841
rect 29089 12832 29101 12835
rect 28960 12804 29101 12832
rect 28960 12792 28966 12804
rect 29089 12801 29101 12804
rect 29135 12801 29147 12835
rect 29089 12795 29147 12801
rect 29365 12835 29423 12841
rect 29365 12801 29377 12835
rect 29411 12801 29423 12835
rect 29365 12795 29423 12801
rect 29638 12792 29644 12844
rect 29696 12792 29702 12844
rect 29822 12792 29828 12844
rect 29880 12792 29886 12844
rect 30558 12841 30564 12844
rect 30552 12795 30564 12841
rect 30558 12792 30564 12795
rect 30616 12792 30622 12844
rect 27890 12764 27896 12776
rect 26016 12736 26188 12764
rect 27540 12736 27896 12764
rect 26016 12724 26022 12736
rect 27540 12696 27568 12736
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 28994 12724 29000 12776
rect 29052 12764 29058 12776
rect 29457 12767 29515 12773
rect 29457 12764 29469 12767
rect 29052 12736 29469 12764
rect 29052 12724 29058 12736
rect 29457 12733 29469 12736
rect 29503 12733 29515 12767
rect 29457 12727 29515 12733
rect 30282 12724 30288 12776
rect 30340 12724 30346 12776
rect 25424 12668 27568 12696
rect 27614 12656 27620 12708
rect 27672 12656 27678 12708
rect 27982 12656 27988 12708
rect 28040 12696 28046 12708
rect 29549 12699 29607 12705
rect 29549 12696 29561 12699
rect 28040 12668 29561 12696
rect 28040 12656 28046 12668
rect 29549 12665 29561 12668
rect 29595 12696 29607 12699
rect 29595 12668 29776 12696
rect 29595 12665 29607 12668
rect 29549 12659 29607 12665
rect 28000 12628 28028 12656
rect 23348 12600 28028 12628
rect 29748 12628 29776 12668
rect 29914 12628 29920 12640
rect 29748 12600 29920 12628
rect 23348 12588 23354 12600
rect 29914 12588 29920 12600
rect 29972 12628 29978 12640
rect 31665 12631 31723 12637
rect 31665 12628 31677 12631
rect 29972 12600 31677 12628
rect 29972 12588 29978 12600
rect 31665 12597 31677 12600
rect 31711 12597 31723 12631
rect 31665 12591 31723 12597
rect 1104 12538 32476 12560
rect 1104 12486 4871 12538
rect 4923 12486 4935 12538
rect 4987 12486 4999 12538
rect 5051 12486 5063 12538
rect 5115 12486 5127 12538
rect 5179 12486 12713 12538
rect 12765 12486 12777 12538
rect 12829 12486 12841 12538
rect 12893 12486 12905 12538
rect 12957 12486 12969 12538
rect 13021 12486 20555 12538
rect 20607 12486 20619 12538
rect 20671 12486 20683 12538
rect 20735 12486 20747 12538
rect 20799 12486 20811 12538
rect 20863 12486 28397 12538
rect 28449 12486 28461 12538
rect 28513 12486 28525 12538
rect 28577 12486 28589 12538
rect 28641 12486 28653 12538
rect 28705 12486 32476 12538
rect 1104 12464 32476 12486
rect 3142 12424 3148 12436
rect 2608 12396 3148 12424
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12257 2559 12291
rect 2501 12251 2559 12257
rect 2516 12152 2544 12251
rect 2608 12229 2636 12396
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 4157 12427 4215 12433
rect 4157 12393 4169 12427
rect 4203 12424 4215 12427
rect 5626 12424 5632 12436
rect 4203 12396 5632 12424
rect 4203 12393 4215 12396
rect 4157 12387 4215 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 7006 12384 7012 12436
rect 7064 12384 7070 12436
rect 9674 12384 9680 12436
rect 9732 12384 9738 12436
rect 11514 12384 11520 12436
rect 11572 12384 11578 12436
rect 13538 12384 13544 12436
rect 13596 12384 13602 12436
rect 13722 12384 13728 12436
rect 13780 12384 13786 12436
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 15436 12396 15485 12424
rect 15436 12384 15442 12396
rect 15473 12393 15485 12396
rect 15519 12393 15531 12427
rect 15473 12387 15531 12393
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 15746 12424 15752 12436
rect 15703 12396 15752 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 16482 12424 16488 12436
rect 15896 12396 16488 12424
rect 15896 12384 15902 12396
rect 16482 12384 16488 12396
rect 16540 12424 16546 12436
rect 17126 12424 17132 12436
rect 16540 12396 17132 12424
rect 16540 12384 16546 12396
rect 17126 12384 17132 12396
rect 17184 12424 17190 12436
rect 17184 12396 21220 12424
rect 17184 12384 17190 12396
rect 2961 12359 3019 12365
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 3326 12356 3332 12368
rect 3007 12328 3332 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 14274 12316 14280 12368
rect 14332 12316 14338 12368
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 15562 12356 15568 12368
rect 15252 12328 15568 12356
rect 15252 12316 15258 12328
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 3200 12260 4261 12288
rect 3200 12248 3206 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6362 12288 6368 12300
rect 5592 12260 6368 12288
rect 5592 12248 5598 12260
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12288 9459 12291
rect 9950 12288 9956 12300
rect 9447 12260 9956 12288
rect 9447 12257 9459 12260
rect 9401 12251 9459 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 15470 12288 15476 12300
rect 14568 12260 15476 12288
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6196 12192 7205 12220
rect 3234 12152 3240 12164
rect 2516 12124 3240 12152
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 6196 12093 6224 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 9180 12192 9321 12220
rect 9180 12180 9186 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12220 10195 12223
rect 11146 12220 11152 12232
rect 10183 12192 11152 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 12066 12180 12072 12232
rect 12124 12180 12130 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 13630 12220 13636 12232
rect 12391 12192 13636 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 14568 12229 14596 12260
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 17221 12223 17279 12229
rect 17221 12220 17233 12223
rect 15304 12192 17233 12220
rect 15304 12164 15332 12192
rect 17221 12189 17233 12192
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 19426 12220 19432 12232
rect 18555 12192 19432 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 21192 12229 21220 12396
rect 21542 12384 21548 12436
rect 21600 12384 21606 12436
rect 22005 12427 22063 12433
rect 22005 12393 22017 12427
rect 22051 12424 22063 12427
rect 22830 12424 22836 12436
rect 22051 12396 22836 12424
rect 22051 12393 22063 12396
rect 22005 12387 22063 12393
rect 22830 12384 22836 12396
rect 22888 12384 22894 12436
rect 23198 12384 23204 12436
rect 23256 12384 23262 12436
rect 26234 12384 26240 12436
rect 26292 12424 26298 12436
rect 26329 12427 26387 12433
rect 26329 12424 26341 12427
rect 26292 12396 26341 12424
rect 26292 12384 26298 12396
rect 26329 12393 26341 12396
rect 26375 12393 26387 12427
rect 26329 12387 26387 12393
rect 27706 12384 27712 12436
rect 27764 12384 27770 12436
rect 30558 12384 30564 12436
rect 30616 12424 30622 12436
rect 30745 12427 30803 12433
rect 30745 12424 30757 12427
rect 30616 12396 30757 12424
rect 30616 12384 30622 12396
rect 30745 12393 30757 12396
rect 30791 12393 30803 12427
rect 30745 12387 30803 12393
rect 23290 12356 23296 12368
rect 22066 12328 23296 12356
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 22066 12288 22094 12328
rect 23290 12316 23296 12328
rect 23348 12356 23354 12368
rect 23348 12328 23428 12356
rect 23348 12316 23354 12328
rect 21315 12260 22094 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 22278 12248 22284 12300
rect 22336 12288 22342 12300
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 22336 12260 22477 12288
rect 22336 12248 22342 12260
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22465 12251 22523 12257
rect 22554 12248 22560 12300
rect 22612 12248 22618 12300
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 23400 12229 23428 12328
rect 24670 12316 24676 12368
rect 24728 12356 24734 12368
rect 28353 12359 28411 12365
rect 28353 12356 28365 12359
rect 24728 12328 28365 12356
rect 24728 12316 24734 12328
rect 28353 12325 28365 12328
rect 28399 12325 28411 12359
rect 28353 12319 28411 12325
rect 29822 12316 29828 12368
rect 29880 12356 29886 12368
rect 29880 12328 30144 12356
rect 29880 12316 29886 12328
rect 25498 12248 25504 12300
rect 25556 12288 25562 12300
rect 25556 12260 25820 12288
rect 25556 12248 25562 12260
rect 25792 12232 25820 12260
rect 25958 12248 25964 12300
rect 26016 12248 26022 12300
rect 29454 12288 29460 12300
rect 29104 12260 29460 12288
rect 29104 12232 29132 12260
rect 29454 12248 29460 12260
rect 29512 12248 29518 12300
rect 30006 12248 30012 12300
rect 30064 12248 30070 12300
rect 30116 12297 30144 12328
rect 30101 12291 30159 12297
rect 30101 12257 30113 12291
rect 30147 12257 30159 12291
rect 30101 12251 30159 12257
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 22796 12192 23213 12220
rect 22796 12180 22802 12192
rect 23201 12189 23213 12192
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 6362 12161 6368 12164
rect 6349 12155 6368 12161
rect 6349 12121 6361 12155
rect 6349 12115 6368 12121
rect 6362 12112 6368 12115
rect 6420 12112 6426 12164
rect 6549 12155 6607 12161
rect 6549 12121 6561 12155
rect 6595 12152 6607 12155
rect 6638 12152 6644 12164
rect 6595 12124 6644 12152
rect 6595 12121 6607 12124
rect 6549 12115 6607 12121
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 10410 12161 10416 12164
rect 10404 12115 10416 12161
rect 10410 12112 10416 12115
rect 10468 12112 10474 12164
rect 13357 12155 13415 12161
rect 13357 12121 13369 12155
rect 13403 12152 13415 12155
rect 13446 12152 13452 12164
rect 13403 12124 13452 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 14645 12155 14703 12161
rect 14645 12121 14657 12155
rect 14691 12152 14703 12155
rect 15194 12152 15200 12164
rect 14691 12124 15200 12152
rect 14691 12121 14703 12124
rect 14645 12115 14703 12121
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 15286 12112 15292 12164
rect 15344 12112 15350 12164
rect 17034 12112 17040 12164
rect 17092 12152 17098 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 17092 12124 18061 12152
rect 17092 12112 17098 12124
rect 18049 12121 18061 12124
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 12161 12087 12219 12093
rect 12161 12053 12173 12087
rect 12207 12084 12219 12087
rect 12434 12084 12440 12096
rect 12207 12056 12440 12084
rect 12207 12053 12219 12056
rect 12161 12047 12219 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12526 12044 12532 12096
rect 12584 12044 12590 12096
rect 13567 12087 13625 12093
rect 13567 12053 13579 12087
rect 13613 12084 13625 12087
rect 13906 12084 13912 12096
rect 13613 12056 13912 12084
rect 13613 12053 13625 12056
rect 13567 12047 13625 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 15470 12044 15476 12096
rect 15528 12093 15534 12096
rect 15528 12087 15557 12093
rect 15545 12084 15557 12087
rect 15838 12084 15844 12096
rect 15545 12056 15844 12084
rect 15545 12053 15557 12056
rect 15528 12047 15557 12053
rect 15528 12044 15534 12047
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 17589 12087 17647 12093
rect 17589 12053 17601 12087
rect 17635 12084 17647 12087
rect 17770 12084 17776 12096
rect 17635 12056 17776 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 18248 12084 18276 12180
rect 18417 12155 18475 12161
rect 18417 12121 18429 12155
rect 18463 12152 18475 12155
rect 18598 12152 18604 12164
rect 18463 12124 18604 12152
rect 18463 12121 18475 12124
rect 18417 12115 18475 12121
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 22094 12112 22100 12164
rect 22152 12152 22158 12164
rect 22373 12155 22431 12161
rect 22373 12152 22385 12155
rect 22152 12124 22385 12152
rect 22152 12112 22158 12124
rect 22373 12121 22385 12124
rect 22419 12152 22431 12155
rect 23658 12152 23664 12164
rect 22419 12124 23664 12152
rect 22419 12121 22431 12124
rect 22373 12115 22431 12121
rect 23658 12112 23664 12124
rect 23716 12112 23722 12164
rect 19150 12084 19156 12096
rect 18248 12056 19156 12084
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 22646 12044 22652 12096
rect 22704 12084 22710 12096
rect 24780 12084 24808 12183
rect 24946 12180 24952 12232
rect 25004 12180 25010 12232
rect 25590 12180 25596 12232
rect 25648 12180 25654 12232
rect 25774 12180 25780 12232
rect 25832 12180 25838 12232
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12189 25927 12223
rect 25869 12183 25927 12189
rect 25682 12112 25688 12164
rect 25740 12152 25746 12164
rect 25884 12152 25912 12183
rect 26050 12180 26056 12232
rect 26108 12220 26114 12232
rect 26145 12223 26203 12229
rect 26145 12220 26157 12223
rect 26108 12192 26157 12220
rect 26108 12180 26114 12192
rect 26145 12189 26157 12192
rect 26191 12189 26203 12223
rect 26145 12183 26203 12189
rect 27985 12223 28043 12229
rect 27985 12189 27997 12223
rect 28031 12189 28043 12223
rect 27985 12183 28043 12189
rect 28445 12223 28503 12229
rect 28445 12189 28457 12223
rect 28491 12220 28503 12223
rect 29086 12220 29092 12232
rect 28491 12192 29092 12220
rect 28491 12189 28503 12192
rect 28445 12183 28503 12189
rect 25740 12124 25912 12152
rect 28000 12152 28028 12183
rect 29086 12180 29092 12192
rect 29144 12180 29150 12232
rect 29181 12223 29239 12229
rect 29181 12189 29193 12223
rect 29227 12220 29239 12223
rect 29638 12220 29644 12232
rect 29227 12192 29644 12220
rect 29227 12189 29239 12192
rect 29181 12183 29239 12189
rect 29638 12180 29644 12192
rect 29696 12180 29702 12232
rect 29917 12223 29975 12229
rect 29917 12189 29929 12223
rect 29963 12189 29975 12223
rect 29917 12183 29975 12189
rect 28905 12155 28963 12161
rect 28000 12124 28856 12152
rect 25740 12112 25746 12124
rect 22704 12056 24808 12084
rect 25133 12087 25191 12093
rect 22704 12044 22710 12056
rect 25133 12053 25145 12087
rect 25179 12084 25191 12087
rect 25314 12084 25320 12096
rect 25179 12056 25320 12084
rect 25179 12053 25191 12056
rect 25133 12047 25191 12053
rect 25314 12044 25320 12056
rect 25372 12084 25378 12096
rect 28074 12084 28080 12096
rect 25372 12056 28080 12084
rect 25372 12044 25378 12056
rect 28074 12044 28080 12056
rect 28132 12044 28138 12096
rect 28166 12044 28172 12096
rect 28224 12044 28230 12096
rect 28828 12084 28856 12124
rect 28905 12121 28917 12155
rect 28951 12152 28963 12155
rect 29270 12152 29276 12164
rect 28951 12124 29276 12152
rect 28951 12121 28963 12124
rect 28905 12115 28963 12121
rect 29270 12112 29276 12124
rect 29328 12112 29334 12164
rect 29932 12152 29960 12183
rect 30190 12180 30196 12232
rect 30248 12180 30254 12232
rect 30742 12180 30748 12232
rect 30800 12220 30806 12232
rect 30929 12223 30987 12229
rect 30929 12220 30941 12223
rect 30800 12192 30941 12220
rect 30800 12180 30806 12192
rect 30929 12189 30941 12192
rect 30975 12189 30987 12223
rect 30929 12183 30987 12189
rect 30374 12152 30380 12164
rect 29932 12124 30380 12152
rect 30374 12112 30380 12124
rect 30432 12112 30438 12164
rect 28994 12084 29000 12096
rect 29052 12093 29058 12096
rect 28828 12056 29000 12084
rect 28994 12044 29000 12056
rect 29052 12047 29061 12093
rect 29052 12044 29058 12047
rect 29730 12044 29736 12096
rect 29788 12044 29794 12096
rect 1104 11994 32632 12016
rect 1104 11942 8792 11994
rect 8844 11942 8856 11994
rect 8908 11942 8920 11994
rect 8972 11942 8984 11994
rect 9036 11942 9048 11994
rect 9100 11942 16634 11994
rect 16686 11942 16698 11994
rect 16750 11942 16762 11994
rect 16814 11942 16826 11994
rect 16878 11942 16890 11994
rect 16942 11942 24476 11994
rect 24528 11942 24540 11994
rect 24592 11942 24604 11994
rect 24656 11942 24668 11994
rect 24720 11942 24732 11994
rect 24784 11942 32318 11994
rect 32370 11942 32382 11994
rect 32434 11942 32446 11994
rect 32498 11942 32510 11994
rect 32562 11942 32574 11994
rect 32626 11942 32632 11994
rect 1104 11920 32632 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11880 3111 11883
rect 4062 11880 4068 11892
rect 3099 11852 4068 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 15470 11880 15476 11892
rect 14884 11852 15476 11880
rect 14884 11840 14890 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 16776 11852 18613 11880
rect 2866 11772 2872 11824
rect 2924 11812 2930 11824
rect 7742 11812 7748 11824
rect 2924 11784 7748 11812
rect 2924 11772 2930 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 10904 11815 10962 11821
rect 10904 11781 10916 11815
rect 10950 11812 10962 11815
rect 12526 11812 12532 11824
rect 10950 11784 12532 11812
rect 10950 11781 10962 11784
rect 10904 11775 10962 11781
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 14642 11772 14648 11824
rect 14700 11772 14706 11824
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 15838 11812 15844 11824
rect 15252 11784 15844 11812
rect 15252 11772 15258 11784
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3602 11744 3608 11756
rect 3292 11716 3608 11744
rect 3292 11704 3298 11716
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4873 11747 4931 11753
rect 4873 11744 4885 11747
rect 4764 11716 4885 11744
rect 4764 11704 4770 11716
rect 4873 11713 4885 11716
rect 4919 11713 4931 11747
rect 4873 11707 4931 11713
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7374 11744 7380 11756
rect 6963 11716 7380 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 13630 11704 13636 11756
rect 13688 11704 13694 11756
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14458 11744 14464 11756
rect 14148 11716 14464 11744
rect 14148 11704 14154 11716
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11744 15439 11747
rect 15562 11744 15568 11756
rect 15427 11716 15568 11744
rect 15427 11713 15439 11716
rect 15381 11707 15439 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16776 11744 16804 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 25774 11840 25780 11892
rect 25832 11880 25838 11892
rect 26421 11883 26479 11889
rect 26421 11880 26433 11883
rect 25832 11852 26433 11880
rect 25832 11840 25838 11852
rect 26421 11849 26433 11852
rect 26467 11849 26479 11883
rect 26421 11843 26479 11849
rect 28166 11840 28172 11892
rect 28224 11840 28230 11892
rect 29362 11840 29368 11892
rect 29420 11840 29426 11892
rect 29917 11883 29975 11889
rect 29917 11849 29929 11883
rect 29963 11880 29975 11883
rect 30190 11880 30196 11892
rect 29963 11852 30196 11880
rect 29963 11849 29975 11852
rect 29917 11843 29975 11849
rect 30190 11840 30196 11852
rect 30248 11840 30254 11892
rect 16945 11815 17003 11821
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 17862 11812 17868 11824
rect 16991 11784 17868 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 17862 11772 17868 11784
rect 17920 11812 17926 11824
rect 18141 11815 18199 11821
rect 18141 11812 18153 11815
rect 17920 11784 18153 11812
rect 17920 11772 17926 11784
rect 18141 11781 18153 11784
rect 18187 11781 18199 11815
rect 23658 11812 23664 11824
rect 18141 11775 18199 11781
rect 23584 11784 23664 11812
rect 16347 11716 16804 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16850 11704 16856 11756
rect 16908 11704 16914 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17218 11744 17224 11756
rect 17083 11716 17224 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17770 11704 17776 11756
rect 17828 11704 17834 11756
rect 18782 11704 18788 11756
rect 18840 11704 18846 11756
rect 18966 11704 18972 11756
rect 19024 11744 19030 11756
rect 19061 11747 19119 11753
rect 19061 11744 19073 11747
rect 19024 11716 19073 11744
rect 19024 11704 19030 11716
rect 19061 11713 19073 11716
rect 19107 11713 19119 11747
rect 19061 11707 19119 11713
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 23584 11753 23612 11784
rect 23658 11772 23664 11784
rect 23716 11812 23722 11824
rect 25682 11812 25688 11824
rect 23716 11784 25688 11812
rect 23716 11772 23722 11784
rect 25682 11772 25688 11784
rect 25740 11772 25746 11824
rect 25958 11772 25964 11824
rect 26016 11812 26022 11824
rect 29730 11812 29736 11824
rect 26016 11784 27200 11812
rect 26016 11772 26022 11784
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 22244 11716 22385 11744
rect 22244 11704 22250 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11744 23811 11747
rect 23934 11744 23940 11756
rect 23799 11716 23940 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 27172 11753 27200 11784
rect 28736 11784 29736 11812
rect 26513 11747 26571 11753
rect 26513 11713 26525 11747
rect 26559 11713 26571 11747
rect 26513 11707 26571 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11744 27215 11747
rect 27614 11744 27620 11756
rect 27203 11716 27620 11744
rect 27203 11713 27215 11716
rect 27157 11707 27215 11713
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 2648 11648 3433 11676
rect 2648 11636 2654 11648
rect 3421 11645 3433 11648
rect 3467 11676 3479 11679
rect 4430 11676 4436 11688
rect 3467 11648 4436 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 5776 11648 7021 11676
rect 5776 11636 5782 11648
rect 7009 11645 7021 11648
rect 7055 11676 7067 11679
rect 10134 11676 10140 11688
rect 7055 11648 10140 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 15109 11679 15167 11685
rect 15109 11676 15121 11679
rect 14608 11648 15121 11676
rect 14608 11636 14614 11648
rect 15109 11645 15121 11648
rect 15155 11676 15167 11679
rect 15289 11679 15347 11685
rect 15155 11648 15240 11676
rect 15155 11645 15167 11648
rect 15109 11639 15167 11645
rect 15212 11608 15240 11648
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 15746 11676 15752 11688
rect 15335 11648 15752 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 17402 11676 17408 11688
rect 16255 11648 17408 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11645 17739 11679
rect 17681 11639 17739 11645
rect 16114 11608 16120 11620
rect 15212 11580 16120 11608
rect 16114 11568 16120 11580
rect 16172 11568 16178 11620
rect 17497 11611 17555 11617
rect 17497 11608 17509 11611
rect 16316 11580 17509 11608
rect 5994 11500 6000 11552
rect 6052 11500 6058 11552
rect 6549 11543 6607 11549
rect 6549 11509 6561 11543
rect 6595 11540 6607 11543
rect 6638 11540 6644 11552
rect 6595 11512 6644 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 7800 11512 9781 11540
rect 7800 11500 7806 11512
rect 9769 11509 9781 11512
rect 9815 11540 9827 11543
rect 12434 11540 12440 11552
rect 9815 11512 12440 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13320 11512 13461 11540
rect 13320 11500 13326 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 14369 11543 14427 11549
rect 14369 11509 14381 11543
rect 14415 11540 14427 11543
rect 14642 11540 14648 11552
rect 14415 11512 14648 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15194 11500 15200 11552
rect 15252 11500 15258 11552
rect 15930 11500 15936 11552
rect 15988 11500 15994 11552
rect 16316 11549 16344 11580
rect 17497 11577 17509 11580
rect 17543 11577 17555 11611
rect 17497 11571 17555 11577
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 17126 11540 17132 11552
rect 16908 11512 17132 11540
rect 16908 11500 16914 11512
rect 17126 11500 17132 11512
rect 17184 11540 17190 11552
rect 17696 11540 17724 11639
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 22465 11679 22523 11685
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 23842 11676 23848 11688
rect 22511 11648 23848 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18892 11608 18920 11639
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 26528 11676 26556 11707
rect 27614 11704 27620 11716
rect 27672 11704 27678 11756
rect 27890 11704 27896 11756
rect 27948 11704 27954 11756
rect 27982 11704 27988 11756
rect 28040 11704 28046 11756
rect 28074 11704 28080 11756
rect 28132 11744 28138 11756
rect 28736 11753 28764 11784
rect 29730 11772 29736 11784
rect 29788 11772 29794 11824
rect 28721 11747 28779 11753
rect 28132 11716 28672 11744
rect 28132 11704 28138 11716
rect 27433 11679 27491 11685
rect 26528 11648 27292 11676
rect 18012 11580 18920 11608
rect 22005 11611 22063 11617
rect 18012 11568 18018 11580
rect 22005 11577 22017 11611
rect 22051 11608 22063 11611
rect 22554 11608 22560 11620
rect 22051 11580 22560 11608
rect 22051 11577 22063 11580
rect 22005 11571 22063 11577
rect 22554 11568 22560 11580
rect 22612 11568 22618 11620
rect 27264 11617 27292 11648
rect 27433 11645 27445 11679
rect 27479 11676 27491 11679
rect 27522 11676 27528 11688
rect 27479 11648 27528 11676
rect 27479 11645 27491 11648
rect 27433 11639 27491 11645
rect 27522 11636 27528 11648
rect 27580 11636 27586 11688
rect 28169 11679 28227 11685
rect 28169 11645 28181 11679
rect 28215 11645 28227 11679
rect 28644 11676 28672 11716
rect 28721 11713 28733 11747
rect 28767 11713 28779 11747
rect 28721 11707 28779 11713
rect 28905 11747 28963 11753
rect 28905 11713 28917 11747
rect 28951 11713 28963 11747
rect 28905 11707 28963 11713
rect 28997 11747 29055 11753
rect 28997 11713 29009 11747
rect 29043 11713 29055 11747
rect 28997 11707 29055 11713
rect 29089 11747 29147 11753
rect 29089 11713 29101 11747
rect 29135 11713 29147 11747
rect 29089 11707 29147 11713
rect 28920 11676 28948 11707
rect 28644 11648 28948 11676
rect 28169 11639 28227 11645
rect 27249 11611 27307 11617
rect 27249 11577 27261 11611
rect 27295 11608 27307 11611
rect 27798 11608 27804 11620
rect 27295 11580 27804 11608
rect 27295 11577 27307 11580
rect 27249 11571 27307 11577
rect 27798 11568 27804 11580
rect 27856 11568 27862 11620
rect 28184 11608 28212 11639
rect 28718 11608 28724 11620
rect 28184 11580 28724 11608
rect 28718 11568 28724 11580
rect 28776 11608 28782 11620
rect 29012 11608 29040 11707
rect 29104 11676 29132 11707
rect 29638 11704 29644 11756
rect 29696 11744 29702 11756
rect 29825 11747 29883 11753
rect 29825 11744 29837 11747
rect 29696 11716 29837 11744
rect 29696 11704 29702 11716
rect 29825 11713 29837 11716
rect 29871 11713 29883 11747
rect 29825 11707 29883 11713
rect 30009 11747 30067 11753
rect 30009 11713 30021 11747
rect 30055 11744 30067 11747
rect 30653 11747 30711 11753
rect 30653 11744 30665 11747
rect 30055 11716 30665 11744
rect 30055 11713 30067 11716
rect 30009 11707 30067 11713
rect 30653 11713 30665 11716
rect 30699 11713 30711 11747
rect 30653 11707 30711 11713
rect 29914 11676 29920 11688
rect 29104 11648 29920 11676
rect 29914 11636 29920 11648
rect 29972 11676 29978 11688
rect 30024 11676 30052 11707
rect 29972 11648 30052 11676
rect 29972 11636 29978 11648
rect 30190 11636 30196 11688
rect 30248 11676 30254 11688
rect 30561 11679 30619 11685
rect 30561 11676 30573 11679
rect 30248 11648 30573 11676
rect 30248 11636 30254 11648
rect 30561 11645 30573 11648
rect 30607 11645 30619 11679
rect 30561 11639 30619 11645
rect 29086 11608 29092 11620
rect 28776 11580 29092 11608
rect 28776 11568 28782 11580
rect 29086 11568 29092 11580
rect 29144 11568 29150 11620
rect 17184 11512 17724 11540
rect 17184 11500 17190 11512
rect 19058 11500 19064 11552
rect 19116 11500 19122 11552
rect 22738 11500 22744 11552
rect 22796 11540 22802 11552
rect 23661 11543 23719 11549
rect 23661 11540 23673 11543
rect 22796 11512 23673 11540
rect 22796 11500 22802 11512
rect 23661 11509 23673 11512
rect 23707 11509 23719 11543
rect 23661 11503 23719 11509
rect 27338 11500 27344 11552
rect 27396 11500 27402 11552
rect 30929 11543 30987 11549
rect 30929 11509 30941 11543
rect 30975 11540 30987 11543
rect 31018 11540 31024 11552
rect 30975 11512 31024 11540
rect 30975 11509 30987 11512
rect 30929 11503 30987 11509
rect 31018 11500 31024 11512
rect 31076 11500 31082 11552
rect 1104 11450 32476 11472
rect 1104 11398 4871 11450
rect 4923 11398 4935 11450
rect 4987 11398 4999 11450
rect 5051 11398 5063 11450
rect 5115 11398 5127 11450
rect 5179 11398 12713 11450
rect 12765 11398 12777 11450
rect 12829 11398 12841 11450
rect 12893 11398 12905 11450
rect 12957 11398 12969 11450
rect 13021 11398 20555 11450
rect 20607 11398 20619 11450
rect 20671 11398 20683 11450
rect 20735 11398 20747 11450
rect 20799 11398 20811 11450
rect 20863 11398 28397 11450
rect 28449 11398 28461 11450
rect 28513 11398 28525 11450
rect 28577 11398 28589 11450
rect 28641 11398 28653 11450
rect 28705 11398 32476 11450
rect 1104 11376 32476 11398
rect 2976 11308 4660 11336
rect 2976 11209 3004 11308
rect 4249 11271 4307 11277
rect 4249 11237 4261 11271
rect 4295 11237 4307 11271
rect 4632 11268 4660 11308
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 4893 11339 4951 11345
rect 4893 11336 4905 11339
rect 4764 11308 4905 11336
rect 4764 11296 4770 11308
rect 4893 11305 4905 11308
rect 4939 11305 4951 11339
rect 4893 11299 4951 11305
rect 5721 11339 5779 11345
rect 5721 11305 5733 11339
rect 5767 11336 5779 11339
rect 5994 11336 6000 11348
rect 5767 11308 6000 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 5736 11268 5764 11299
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 9766 11296 9772 11348
rect 9824 11296 9830 11348
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 15286 11336 15292 11348
rect 12406 11308 15292 11336
rect 4632 11240 5764 11268
rect 6549 11271 6607 11277
rect 4249 11231 4307 11237
rect 6549 11237 6561 11271
rect 6595 11268 6607 11271
rect 6638 11268 6644 11280
rect 6595 11240 6644 11268
rect 6595 11237 6607 11240
rect 6549 11231 6607 11237
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4264 11132 4292 11231
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 6917 11271 6975 11277
rect 6917 11237 6929 11271
rect 6963 11268 6975 11271
rect 12406 11268 12434 11308
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16853 11339 16911 11345
rect 16853 11305 16865 11339
rect 16899 11336 16911 11339
rect 17034 11336 17040 11348
rect 16899 11308 17040 11336
rect 16899 11305 16911 11308
rect 16853 11299 16911 11305
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 17460 11308 17509 11336
rect 17460 11296 17466 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 19426 11296 19432 11348
rect 19484 11296 19490 11348
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 23934 11336 23940 11348
rect 22428 11308 23940 11336
rect 22428 11296 22434 11308
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 25130 11296 25136 11348
rect 25188 11296 25194 11348
rect 25866 11296 25872 11348
rect 25924 11336 25930 11348
rect 29825 11339 29883 11345
rect 29825 11336 29837 11339
rect 25924 11308 29837 11336
rect 25924 11296 25930 11308
rect 29825 11305 29837 11308
rect 29871 11336 29883 11339
rect 29871 11308 30052 11336
rect 29871 11305 29883 11308
rect 29825 11299 29883 11305
rect 6963 11240 12434 11268
rect 6963 11237 6975 11240
rect 6917 11231 6975 11237
rect 13630 11228 13636 11280
rect 13688 11268 13694 11280
rect 16669 11271 16727 11277
rect 16669 11268 16681 11271
rect 13688 11240 16681 11268
rect 13688 11228 13694 11240
rect 16669 11237 16681 11240
rect 16715 11237 16727 11271
rect 16669 11231 16727 11237
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 17828 11240 18184 11268
rect 17828 11228 17834 11240
rect 5626 11200 5632 11212
rect 5092 11172 5632 11200
rect 5092 11141 5120 11172
rect 5626 11160 5632 11172
rect 5684 11200 5690 11212
rect 15473 11203 15531 11209
rect 5684 11172 7788 11200
rect 5684 11160 5690 11172
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4264 11104 4905 11132
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 6052 11104 6469 11132
rect 6052 11092 6058 11104
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7558 11132 7564 11144
rect 6779 11104 7564 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 5705 11067 5763 11073
rect 4295 11036 5580 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 2501 10999 2559 11005
rect 2501 10965 2513 10999
rect 2547 10996 2559 10999
rect 2590 10996 2596 11008
rect 2547 10968 2596 10996
rect 2547 10965 2559 10968
rect 2501 10959 2559 10965
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 5552 11005 5580 11036
rect 5705 11033 5717 11067
rect 5751 11064 5763 11067
rect 5810 11064 5816 11076
rect 5751 11036 5816 11064
rect 5751 11033 5763 11036
rect 5705 11027 5763 11033
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 5902 11024 5908 11076
rect 5960 11024 5966 11076
rect 6086 11024 6092 11076
rect 6144 11064 6150 11076
rect 6656 11064 6684 11095
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 7760 11141 7788 11172
rect 8312 11172 10640 11200
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11132 7803 11135
rect 8110 11132 8116 11144
rect 7791 11104 8116 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 6822 11064 6828 11076
rect 6144 11036 6828 11064
rect 6144 11024 6150 11036
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7377 11067 7435 11073
rect 7377 11064 7389 11067
rect 7248 11036 7389 11064
rect 7248 11024 7254 11036
rect 7377 11033 7389 11036
rect 7423 11064 7435 11067
rect 8312 11064 8340 11172
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 7423 11036 8340 11064
rect 8404 11064 8432 11095
rect 9674 11092 9680 11144
rect 9732 11092 9738 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10612 11141 10640 11172
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15654 11200 15660 11212
rect 15519 11172 15660 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 18046 11200 18052 11212
rect 17696 11172 18052 11200
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 10284 11104 10425 11132
rect 10284 11092 10290 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 11054 11132 11060 11144
rect 10643 11104 11060 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 11054 11092 11060 11104
rect 11112 11132 11118 11144
rect 11882 11132 11888 11144
rect 11112 11104 11888 11132
rect 11112 11092 11118 11104
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14366 11132 14372 11144
rect 14323 11104 14372 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 14826 11132 14832 11144
rect 14599 11104 14832 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 17696 11141 17724 11172
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 18156 11209 18184 11240
rect 19058 11228 19064 11280
rect 19116 11268 19122 11280
rect 20165 11271 20223 11277
rect 20165 11268 20177 11271
rect 19116 11240 20177 11268
rect 19116 11228 19122 11240
rect 20165 11237 20177 11240
rect 20211 11268 20223 11271
rect 22557 11271 22615 11277
rect 22557 11268 22569 11271
rect 20211 11240 22569 11268
rect 20211 11237 20223 11240
rect 20165 11231 20223 11237
rect 22557 11237 22569 11240
rect 22603 11237 22615 11271
rect 23750 11268 23756 11280
rect 22557 11231 22615 11237
rect 22756 11240 23756 11268
rect 18141 11203 18199 11209
rect 18141 11169 18153 11203
rect 18187 11200 18199 11203
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 18187 11172 19717 11200
rect 18187 11169 18199 11172
rect 18141 11163 18199 11169
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 20717 11203 20775 11209
rect 20717 11200 20729 11203
rect 19705 11163 19763 11169
rect 20180 11172 20729 11200
rect 17681 11135 17739 11141
rect 17681 11132 17693 11135
rect 15620 11104 17693 11132
rect 15620 11092 15626 11104
rect 17681 11101 17693 11104
rect 17727 11101 17739 11135
rect 17681 11095 17739 11101
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11132 17831 11135
rect 17862 11132 17868 11144
rect 17819 11104 17868 11132
rect 17819 11101 17831 11104
rect 17773 11095 17831 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 20180 11076 20208 11172
rect 20717 11169 20729 11172
rect 20763 11169 20775 11203
rect 20717 11163 20775 11169
rect 20993 11203 21051 11209
rect 20993 11169 21005 11203
rect 21039 11169 21051 11203
rect 22756 11200 22784 11240
rect 23750 11228 23756 11240
rect 23808 11268 23814 11280
rect 26789 11271 26847 11277
rect 23808 11240 24808 11268
rect 23808 11228 23814 11240
rect 23569 11203 23627 11209
rect 23569 11200 23581 11203
rect 20993 11163 21051 11169
rect 21100 11172 22784 11200
rect 22848 11172 23581 11200
rect 20254 11092 20260 11144
rect 20312 11132 20318 11144
rect 21008 11132 21036 11163
rect 21100 11141 21128 11172
rect 20312 11104 21036 11132
rect 21085 11135 21143 11141
rect 20312 11092 20318 11104
rect 21085 11101 21097 11135
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 22848 11141 22876 11172
rect 23569 11169 23581 11172
rect 23615 11169 23627 11203
rect 23569 11163 23627 11169
rect 23658 11160 23664 11212
rect 23716 11160 23722 11212
rect 24673 11203 24731 11209
rect 24673 11169 24685 11203
rect 24719 11169 24731 11203
rect 24673 11163 24731 11169
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11101 22891 11135
rect 22833 11095 22891 11101
rect 23106 11092 23112 11144
rect 23164 11092 23170 11144
rect 23676 11132 23704 11160
rect 23753 11135 23811 11141
rect 23753 11132 23765 11135
rect 23676 11104 23765 11132
rect 23753 11101 23765 11104
rect 23799 11101 23811 11135
rect 23753 11095 23811 11101
rect 23934 11092 23940 11144
rect 23992 11092 23998 11144
rect 10042 11064 10048 11076
rect 8404 11036 10048 11064
rect 7423 11033 7435 11036
rect 7377 11027 7435 11033
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 14737 11067 14795 11073
rect 14737 11033 14749 11067
rect 14783 11064 14795 11067
rect 15470 11064 15476 11076
rect 14783 11036 15476 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 15930 11024 15936 11076
rect 15988 11064 15994 11076
rect 16821 11067 16879 11073
rect 16821 11064 16833 11067
rect 15988 11036 16833 11064
rect 15988 11024 15994 11036
rect 16821 11033 16833 11036
rect 16867 11033 16879 11067
rect 16821 11027 16879 11033
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 17037 11067 17095 11073
rect 17037 11064 17049 11067
rect 17000 11036 17049 11064
rect 17000 11024 17006 11036
rect 17037 11033 17049 11036
rect 17083 11033 17095 11067
rect 17037 11027 17095 11033
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 3476 10968 4077 10996
rect 3476 10956 3482 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 4065 10959 4123 10965
rect 5537 10999 5595 11005
rect 5537 10965 5549 10999
rect 5583 10965 5595 10999
rect 5537 10959 5595 10965
rect 8570 10956 8576 11008
rect 8628 10956 8634 11008
rect 14369 10999 14427 11005
rect 14369 10965 14381 10999
rect 14415 10996 14427 10999
rect 14550 10996 14556 11008
rect 14415 10968 14556 10996
rect 14415 10965 14427 10968
rect 14369 10959 14427 10965
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 15746 10956 15752 11008
rect 15804 10956 15810 11008
rect 17052 10996 17080 11027
rect 17126 11024 17132 11076
rect 17184 11064 17190 11076
rect 18049 11067 18107 11073
rect 18049 11064 18061 11067
rect 17184 11036 18061 11064
rect 17184 11024 17190 11036
rect 18049 11033 18061 11036
rect 18095 11033 18107 11067
rect 18049 11027 18107 11033
rect 20162 11024 20168 11076
rect 20220 11024 20226 11076
rect 22925 11067 22983 11073
rect 22925 11033 22937 11067
rect 22971 11064 22983 11067
rect 23658 11064 23664 11076
rect 22971 11036 23664 11064
rect 22971 11033 22983 11036
rect 22925 11027 22983 11033
rect 23658 11024 23664 11036
rect 23716 11024 23722 11076
rect 24688 11064 24716 11163
rect 24780 11141 24808 11240
rect 26789 11237 26801 11271
rect 26835 11268 26847 11271
rect 27430 11268 27436 11280
rect 26835 11240 27436 11268
rect 26835 11237 26847 11240
rect 26789 11231 26847 11237
rect 27430 11228 27436 11240
rect 27488 11228 27494 11280
rect 28169 11271 28227 11277
rect 28169 11237 28181 11271
rect 28215 11268 28227 11271
rect 29089 11271 29147 11277
rect 29089 11268 29101 11271
rect 28215 11240 29101 11268
rect 28215 11237 28227 11240
rect 28169 11231 28227 11237
rect 29089 11237 29101 11240
rect 29135 11268 29147 11271
rect 30024 11268 30052 11308
rect 30190 11296 30196 11348
rect 30248 11296 30254 11348
rect 30742 11296 30748 11348
rect 30800 11296 30806 11348
rect 30926 11296 30932 11348
rect 30984 11296 30990 11348
rect 31938 11268 31944 11280
rect 29135 11240 29960 11268
rect 30024 11240 31944 11268
rect 29135 11237 29147 11240
rect 29089 11231 29147 11237
rect 27614 11160 27620 11212
rect 27672 11160 27678 11212
rect 28994 11160 29000 11212
rect 29052 11200 29058 11212
rect 29052 11172 29776 11200
rect 29052 11160 29058 11172
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 25774 11092 25780 11144
rect 25832 11092 25838 11144
rect 25866 11092 25872 11144
rect 25924 11092 25930 11144
rect 26513 11135 26571 11141
rect 26513 11101 26525 11135
rect 26559 11132 26571 11135
rect 27798 11132 27804 11144
rect 26559 11104 27804 11132
rect 26559 11101 26571 11104
rect 26513 11095 26571 11101
rect 27798 11092 27804 11104
rect 27856 11092 27862 11144
rect 27982 11092 27988 11144
rect 28040 11092 28046 11144
rect 28905 11135 28963 11141
rect 28905 11101 28917 11135
rect 28951 11101 28963 11135
rect 28905 11095 28963 11101
rect 26789 11067 26847 11073
rect 26789 11064 26801 11067
rect 24688 11036 24900 11064
rect 17402 10996 17408 11008
rect 17052 10968 17408 10996
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 19610 10956 19616 11008
rect 19668 10956 19674 11008
rect 24872 10996 24900 11036
rect 25976 11036 26801 11064
rect 24946 10996 24952 11008
rect 24872 10968 24952 10996
rect 24946 10956 24952 10968
rect 25004 10996 25010 11008
rect 25976 10996 26004 11036
rect 26789 11033 26801 11036
rect 26835 11064 26847 11067
rect 27522 11064 27528 11076
rect 26835 11036 27528 11064
rect 26835 11033 26847 11036
rect 26789 11027 26847 11033
rect 27522 11024 27528 11036
rect 27580 11064 27586 11076
rect 27893 11067 27951 11073
rect 27893 11064 27905 11067
rect 27580 11036 27905 11064
rect 27580 11024 27586 11036
rect 27893 11033 27905 11036
rect 27939 11064 27951 11067
rect 28258 11064 28264 11076
rect 27939 11036 28264 11064
rect 27939 11033 27951 11036
rect 27893 11027 27951 11033
rect 28258 11024 28264 11036
rect 28316 11024 28322 11076
rect 28920 11064 28948 11095
rect 29178 11092 29184 11144
rect 29236 11092 29242 11144
rect 29748 11141 29776 11172
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 29270 11064 29276 11076
rect 28920 11036 29276 11064
rect 29270 11024 29276 11036
rect 29328 11024 29334 11076
rect 29932 11064 29960 11240
rect 31938 11228 31944 11240
rect 31996 11228 32002 11280
rect 31018 11160 31024 11212
rect 31076 11160 31082 11212
rect 31294 11092 31300 11144
rect 31352 11092 31358 11144
rect 30374 11064 30380 11076
rect 29932 11036 30380 11064
rect 30374 11024 30380 11036
rect 30432 11064 30438 11076
rect 30742 11064 30748 11076
rect 30432 11036 30748 11064
rect 30432 11024 30438 11036
rect 30742 11024 30748 11036
rect 30800 11024 30806 11076
rect 25004 10968 26004 10996
rect 25004 10956 25010 10968
rect 26050 10956 26056 11008
rect 26108 10956 26114 11008
rect 26605 10999 26663 11005
rect 26605 10965 26617 10999
rect 26651 10996 26663 10999
rect 27614 10996 27620 11008
rect 26651 10968 27620 10996
rect 26651 10965 26663 10968
rect 26605 10959 26663 10965
rect 27614 10956 27620 10968
rect 27672 10956 27678 11008
rect 27798 10956 27804 11008
rect 27856 10956 27862 11008
rect 28718 10956 28724 11008
rect 28776 10956 28782 11008
rect 1104 10906 32632 10928
rect 1104 10854 8792 10906
rect 8844 10854 8856 10906
rect 8908 10854 8920 10906
rect 8972 10854 8984 10906
rect 9036 10854 9048 10906
rect 9100 10854 16634 10906
rect 16686 10854 16698 10906
rect 16750 10854 16762 10906
rect 16814 10854 16826 10906
rect 16878 10854 16890 10906
rect 16942 10854 24476 10906
rect 24528 10854 24540 10906
rect 24592 10854 24604 10906
rect 24656 10854 24668 10906
rect 24720 10854 24732 10906
rect 24784 10854 32318 10906
rect 32370 10854 32382 10906
rect 32434 10854 32446 10906
rect 32498 10854 32510 10906
rect 32562 10854 32574 10906
rect 32626 10854 32632 10906
rect 1104 10832 32632 10854
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10792 2651 10795
rect 3418 10792 3424 10804
rect 2639 10764 3424 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 3605 10795 3663 10801
rect 3605 10761 3617 10795
rect 3651 10792 3663 10795
rect 3970 10792 3976 10804
rect 3651 10764 3976 10792
rect 3651 10761 3663 10764
rect 3605 10755 3663 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 10042 10752 10048 10804
rect 10100 10752 10106 10804
rect 15286 10792 15292 10804
rect 15212 10764 15292 10792
rect 9585 10727 9643 10733
rect 2746 10696 3464 10724
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2746 10656 2774 10696
rect 2372 10628 2774 10656
rect 2372 10616 2378 10628
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3436 10665 3464 10696
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 9631 10696 13001 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 12989 10693 13001 10696
rect 13035 10724 13047 10727
rect 13078 10724 13084 10736
rect 13035 10696 13084 10724
rect 13035 10693 13047 10696
rect 12989 10687 13047 10693
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 14458 10684 14464 10736
rect 14516 10724 14522 10736
rect 14734 10724 14740 10736
rect 14516 10696 14740 10724
rect 14516 10684 14522 10696
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5718 10656 5724 10668
rect 5399 10628 5724 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6454 10656 6460 10668
rect 5859 10628 6460 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 10226 10616 10232 10668
rect 10284 10616 10290 10668
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 15212 10665 15240 10764
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15654 10792 15660 10804
rect 15488 10764 15660 10792
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15488 10665 15516 10764
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 15838 10752 15844 10804
rect 15896 10752 15902 10804
rect 17405 10795 17463 10801
rect 17405 10761 17417 10795
rect 17451 10792 17463 10795
rect 17954 10792 17960 10804
rect 17451 10764 17960 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 18141 10795 18199 10801
rect 18141 10761 18153 10795
rect 18187 10792 18199 10795
rect 18966 10792 18972 10804
rect 18187 10764 18972 10792
rect 18187 10761 18199 10764
rect 18141 10755 18199 10761
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19076 10764 19809 10792
rect 17218 10724 17224 10736
rect 15580 10696 17224 10724
rect 15580 10665 15608 10696
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15436 10628 15485 10656
rect 15436 10616 15442 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 2590 10548 2596 10600
rect 2648 10588 2654 10600
rect 3329 10591 3387 10597
rect 2648 10560 3004 10588
rect 2648 10548 2654 10560
rect 2409 10523 2467 10529
rect 2409 10489 2421 10523
rect 2455 10520 2467 10523
rect 2682 10520 2688 10532
rect 2455 10492 2688 10520
rect 2455 10489 2467 10492
rect 2409 10483 2467 10489
rect 2682 10480 2688 10492
rect 2740 10520 2746 10532
rect 2976 10520 3004 10560
rect 3329 10557 3341 10591
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 3237 10523 3295 10529
rect 3237 10520 3249 10523
rect 2740 10480 2774 10520
rect 2976 10492 3249 10520
rect 3237 10489 3249 10492
rect 3283 10489 3295 10523
rect 3237 10483 3295 10489
rect 2746 10452 2774 10480
rect 3344 10452 3372 10551
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 9824 10560 10425 10588
rect 9824 10548 9830 10560
rect 10413 10557 10425 10560
rect 10459 10588 10471 10591
rect 10459 10560 12434 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 8662 10520 8668 10532
rect 3476 10492 8668 10520
rect 3476 10480 3482 10492
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 12406 10520 12434 10560
rect 13722 10548 13728 10600
rect 13780 10588 13786 10600
rect 15580 10588 15608 10619
rect 15654 10616 15660 10668
rect 15712 10616 15718 10668
rect 15746 10616 15752 10668
rect 15804 10656 15810 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 15804 10628 17049 10656
rect 15804 10616 15810 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 13780 10560 15608 10588
rect 13780 10548 13786 10560
rect 13630 10520 13636 10532
rect 12406 10492 13636 10520
rect 13630 10480 13636 10492
rect 13688 10480 13694 10532
rect 17052 10520 17080 10619
rect 18322 10616 18328 10668
rect 18380 10616 18386 10668
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 17310 10588 17316 10600
rect 17175 10560 17316 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 18230 10548 18236 10600
rect 18288 10588 18294 10600
rect 18432 10588 18460 10619
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18564 10628 18613 10656
rect 18564 10616 18570 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10656 18751 10659
rect 19076 10656 19104 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 23474 10792 23480 10804
rect 22060 10764 23480 10792
rect 22060 10752 22066 10764
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 25590 10752 25596 10804
rect 25648 10752 25654 10804
rect 27982 10752 27988 10804
rect 28040 10792 28046 10804
rect 28810 10792 28816 10804
rect 28040 10764 28816 10792
rect 28040 10752 28046 10764
rect 28810 10752 28816 10764
rect 28868 10792 28874 10804
rect 31110 10792 31116 10804
rect 28868 10764 31116 10792
rect 28868 10752 28874 10764
rect 19150 10684 19156 10736
rect 19208 10684 19214 10736
rect 19260 10696 22692 10724
rect 18739 10628 19104 10656
rect 18739 10625 18751 10628
rect 18693 10619 18751 10625
rect 18288 10560 18460 10588
rect 18288 10548 18294 10560
rect 18782 10520 18788 10532
rect 17052 10492 18788 10520
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 2746 10424 3372 10452
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 5258 10452 5264 10464
rect 5215 10424 5264 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6822 10452 6828 10464
rect 6043 10424 6828 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 9674 10452 9680 10464
rect 8343 10424 9680 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10452 11759 10455
rect 11790 10452 11796 10464
rect 11747 10424 11796 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 19260 10452 19288 10696
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 19794 10656 19800 10668
rect 19659 10628 19800 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 19794 10616 19800 10628
rect 19852 10616 19858 10668
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19392 10560 19441 10588
rect 19392 10548 19398 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 19518 10548 19524 10600
rect 19576 10588 19582 10600
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 19576 10560 20545 10588
rect 19576 10548 19582 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 20640 10588 20668 10619
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 22186 10616 22192 10668
rect 22244 10616 22250 10668
rect 22296 10665 22324 10696
rect 22281 10659 22339 10665
rect 22281 10625 22293 10659
rect 22327 10625 22339 10659
rect 22281 10619 22339 10625
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10656 22431 10659
rect 22554 10656 22560 10668
rect 22419 10628 22560 10656
rect 22419 10625 22431 10628
rect 22373 10619 22431 10625
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 22664 10656 22692 10696
rect 23382 10684 23388 10736
rect 23440 10684 23446 10736
rect 26510 10724 26516 10736
rect 23492 10696 26516 10724
rect 23290 10656 23296 10668
rect 22664 10628 23296 10656
rect 23290 10616 23296 10628
rect 23348 10656 23354 10668
rect 23492 10656 23520 10696
rect 26510 10684 26516 10696
rect 26568 10684 26574 10736
rect 26602 10684 26608 10736
rect 26660 10724 26666 10736
rect 29178 10724 29184 10736
rect 26660 10696 29184 10724
rect 26660 10684 26666 10696
rect 29178 10684 29184 10696
rect 29236 10684 29242 10736
rect 23348 10628 23520 10656
rect 25961 10659 26019 10665
rect 23348 10616 23354 10628
rect 25961 10625 25973 10659
rect 26007 10625 26019 10659
rect 25961 10619 26019 10625
rect 22462 10588 22468 10600
rect 20640 10560 22468 10588
rect 20533 10551 20591 10557
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 21910 10480 21916 10532
rect 21968 10520 21974 10532
rect 25976 10520 26004 10619
rect 27338 10616 27344 10668
rect 27396 10656 27402 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27396 10628 27537 10656
rect 27396 10616 27402 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 27709 10659 27767 10665
rect 27709 10625 27721 10659
rect 27755 10656 27767 10659
rect 27890 10656 27896 10668
rect 27755 10628 27896 10656
rect 27755 10625 27767 10628
rect 27709 10619 27767 10625
rect 27890 10616 27896 10628
rect 27948 10616 27954 10668
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 28902 10616 28908 10668
rect 28960 10616 28966 10668
rect 29196 10656 29224 10684
rect 29730 10656 29736 10668
rect 29196 10628 29736 10656
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 29840 10665 29868 10764
rect 31110 10752 31116 10764
rect 31168 10792 31174 10804
rect 31297 10795 31355 10801
rect 31297 10792 31309 10795
rect 31168 10764 31309 10792
rect 31168 10752 31174 10764
rect 31297 10761 31309 10764
rect 31343 10761 31355 10795
rect 31297 10755 31355 10761
rect 30098 10684 30104 10736
rect 30156 10724 30162 10736
rect 30469 10727 30527 10733
rect 30469 10724 30481 10727
rect 30156 10696 30481 10724
rect 30156 10684 30162 10696
rect 30469 10693 30481 10696
rect 30515 10693 30527 10727
rect 30469 10687 30527 10693
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10625 29883 10659
rect 29825 10619 29883 10625
rect 30006 10616 30012 10668
rect 30064 10616 30070 10668
rect 30653 10659 30711 10665
rect 30653 10656 30665 10659
rect 30116 10628 30665 10656
rect 26053 10591 26111 10597
rect 26053 10557 26065 10591
rect 26099 10588 26111 10591
rect 27982 10588 27988 10600
rect 26099 10560 27988 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 27982 10548 27988 10560
rect 28040 10548 28046 10600
rect 28626 10548 28632 10600
rect 28684 10588 28690 10600
rect 28813 10591 28871 10597
rect 28813 10588 28825 10591
rect 28684 10560 28825 10588
rect 28684 10548 28690 10560
rect 28813 10557 28825 10560
rect 28859 10557 28871 10591
rect 28813 10551 28871 10557
rect 28994 10548 29000 10600
rect 29052 10548 29058 10600
rect 29748 10588 29776 10616
rect 30116 10588 30144 10628
rect 30653 10625 30665 10628
rect 30699 10625 30711 10659
rect 30653 10619 30711 10625
rect 30742 10616 30748 10668
rect 30800 10616 30806 10668
rect 31205 10659 31263 10665
rect 31205 10625 31217 10659
rect 31251 10656 31263 10659
rect 31294 10656 31300 10668
rect 31251 10628 31300 10656
rect 31251 10625 31263 10628
rect 31205 10619 31263 10625
rect 29748 10560 30144 10588
rect 30558 10548 30564 10600
rect 30616 10588 30622 10600
rect 31220 10588 31248 10619
rect 31294 10616 31300 10628
rect 31352 10616 31358 10668
rect 31481 10659 31539 10665
rect 31481 10625 31493 10659
rect 31527 10656 31539 10659
rect 31754 10656 31760 10668
rect 31527 10628 31760 10656
rect 31527 10625 31539 10628
rect 31481 10619 31539 10625
rect 31754 10616 31760 10628
rect 31812 10616 31818 10668
rect 30616 10560 31248 10588
rect 30616 10548 30622 10560
rect 21968 10492 26004 10520
rect 21968 10480 21974 10492
rect 26326 10480 26332 10532
rect 26384 10520 26390 10532
rect 29181 10523 29239 10529
rect 29181 10520 29193 10523
rect 26384 10492 29193 10520
rect 26384 10480 26390 10492
rect 29181 10489 29193 10492
rect 29227 10489 29239 10523
rect 29181 10483 29239 10489
rect 29270 10480 29276 10532
rect 29328 10520 29334 10532
rect 30469 10523 30527 10529
rect 30469 10520 30481 10523
rect 29328 10492 30481 10520
rect 29328 10480 29334 10492
rect 30469 10489 30481 10492
rect 30515 10489 30527 10523
rect 30469 10483 30527 10489
rect 13596 10424 19288 10452
rect 19613 10455 19671 10461
rect 13596 10412 13602 10424
rect 19613 10421 19625 10455
rect 19659 10452 19671 10455
rect 20162 10452 20168 10464
rect 19659 10424 20168 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 20346 10412 20352 10464
rect 20404 10412 20410 10464
rect 22462 10412 22468 10464
rect 22520 10452 22526 10464
rect 22649 10455 22707 10461
rect 22649 10452 22661 10455
rect 22520 10424 22661 10452
rect 22520 10412 22526 10424
rect 22649 10421 22661 10424
rect 22695 10421 22707 10455
rect 22649 10415 22707 10421
rect 24394 10412 24400 10464
rect 24452 10452 24458 10464
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24452 10424 24685 10452
rect 24452 10412 24458 10424
rect 24673 10421 24685 10424
rect 24719 10421 24731 10455
rect 24673 10415 24731 10421
rect 27614 10412 27620 10464
rect 27672 10452 27678 10464
rect 27893 10455 27951 10461
rect 27893 10452 27905 10455
rect 27672 10424 27905 10452
rect 27672 10412 27678 10424
rect 27893 10421 27905 10424
rect 27939 10421 27951 10455
rect 27893 10415 27951 10421
rect 29638 10412 29644 10464
rect 29696 10412 29702 10464
rect 29730 10412 29736 10464
rect 29788 10452 29794 10464
rect 29825 10455 29883 10461
rect 29825 10452 29837 10455
rect 29788 10424 29837 10452
rect 29788 10412 29794 10424
rect 29825 10421 29837 10424
rect 29871 10421 29883 10455
rect 29825 10415 29883 10421
rect 31018 10412 31024 10464
rect 31076 10452 31082 10464
rect 31481 10455 31539 10461
rect 31481 10452 31493 10455
rect 31076 10424 31493 10452
rect 31076 10412 31082 10424
rect 31481 10421 31493 10424
rect 31527 10421 31539 10455
rect 31481 10415 31539 10421
rect 1104 10362 32476 10384
rect 1104 10310 4871 10362
rect 4923 10310 4935 10362
rect 4987 10310 4999 10362
rect 5051 10310 5063 10362
rect 5115 10310 5127 10362
rect 5179 10310 12713 10362
rect 12765 10310 12777 10362
rect 12829 10310 12841 10362
rect 12893 10310 12905 10362
rect 12957 10310 12969 10362
rect 13021 10310 20555 10362
rect 20607 10310 20619 10362
rect 20671 10310 20683 10362
rect 20735 10310 20747 10362
rect 20799 10310 20811 10362
rect 20863 10310 28397 10362
rect 28449 10310 28461 10362
rect 28513 10310 28525 10362
rect 28577 10310 28589 10362
rect 28641 10310 28653 10362
rect 28705 10310 32476 10362
rect 1104 10288 32476 10310
rect 2682 10208 2688 10260
rect 2740 10208 2746 10260
rect 3050 10208 3056 10260
rect 3108 10208 3114 10260
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3510 10248 3516 10260
rect 3191 10220 3516 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3160 10180 3188 10211
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 6144 10220 7941 10248
rect 6144 10208 6150 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10505 10251 10563 10257
rect 10505 10248 10517 10251
rect 10192 10220 10517 10248
rect 10192 10208 10198 10220
rect 10505 10217 10517 10220
rect 10551 10217 10563 10251
rect 10505 10211 10563 10217
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 15286 10248 15292 10260
rect 14323 10220 15292 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 15620 10220 17509 10248
rect 15620 10208 15626 10220
rect 17497 10217 17509 10220
rect 17543 10248 17555 10251
rect 18414 10248 18420 10260
rect 17543 10220 18420 10248
rect 17543 10217 17555 10220
rect 17497 10211 17555 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18693 10251 18751 10257
rect 18693 10248 18705 10251
rect 18656 10220 18705 10248
rect 18656 10208 18662 10220
rect 18693 10217 18705 10220
rect 18739 10248 18751 10251
rect 19518 10248 19524 10260
rect 18739 10220 19524 10248
rect 18739 10217 18751 10220
rect 18693 10211 18751 10217
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 19981 10251 20039 10257
rect 19981 10248 19993 10251
rect 19668 10220 19993 10248
rect 19668 10208 19674 10220
rect 19981 10217 19993 10220
rect 20027 10217 20039 10251
rect 19981 10211 20039 10217
rect 23017 10251 23075 10257
rect 23017 10217 23029 10251
rect 23063 10248 23075 10251
rect 23106 10248 23112 10260
rect 23063 10220 23112 10248
rect 23063 10217 23075 10220
rect 23017 10211 23075 10217
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 23658 10208 23664 10260
rect 23716 10248 23722 10260
rect 23937 10251 23995 10257
rect 23937 10248 23949 10251
rect 23716 10220 23949 10248
rect 23716 10208 23722 10220
rect 23937 10217 23949 10220
rect 23983 10217 23995 10251
rect 23937 10211 23995 10217
rect 27614 10208 27620 10260
rect 27672 10208 27678 10260
rect 31018 10208 31024 10260
rect 31076 10208 31082 10260
rect 31754 10208 31760 10260
rect 31812 10208 31818 10260
rect 2056 10152 3188 10180
rect 3237 10183 3295 10189
rect 2056 10053 2084 10152
rect 3237 10149 3249 10183
rect 3283 10180 3295 10183
rect 3786 10180 3792 10192
rect 3283 10152 3792 10180
rect 3283 10149 3295 10152
rect 3237 10143 3295 10149
rect 3786 10140 3792 10152
rect 3844 10180 3850 10192
rect 4154 10180 4160 10192
rect 3844 10152 4160 10180
rect 3844 10140 3850 10152
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 15105 10183 15163 10189
rect 15105 10149 15117 10183
rect 15151 10180 15163 10183
rect 15654 10180 15660 10192
rect 15151 10152 15660 10180
rect 15151 10149 15163 10152
rect 15105 10143 15163 10149
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 18506 10140 18512 10192
rect 18564 10140 18570 10192
rect 18782 10140 18788 10192
rect 18840 10180 18846 10192
rect 19429 10183 19487 10189
rect 19429 10180 19441 10183
rect 18840 10152 19441 10180
rect 18840 10140 18846 10152
rect 19429 10149 19441 10152
rect 19475 10149 19487 10183
rect 19429 10143 19487 10149
rect 23198 10140 23204 10192
rect 23256 10180 23262 10192
rect 26786 10180 26792 10192
rect 23256 10152 26792 10180
rect 23256 10140 23262 10152
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10112 14703 10115
rect 15010 10112 15016 10124
rect 14691 10084 15016 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2271 10016 2973 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2961 10013 2973 10016
rect 3007 10044 3019 10047
rect 3326 10044 3332 10056
rect 3007 10016 3332 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3602 10044 3608 10056
rect 3467 10016 3608 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3602 10004 3608 10016
rect 3660 10044 3666 10056
rect 3878 10044 3884 10056
rect 3660 10016 3884 10044
rect 3660 10004 3666 10016
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 6546 10044 6552 10056
rect 4672 10016 6552 10044
rect 4672 10004 4678 10016
rect 6546 10004 6552 10016
rect 6604 10044 6610 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 6604 10016 9137 10044
rect 6604 10004 6610 10016
rect 9125 10013 9137 10016
rect 9171 10044 9183 10047
rect 9674 10044 9680 10056
rect 9171 10016 9680 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9674 10004 9680 10016
rect 9732 10044 9738 10056
rect 11057 10047 11115 10053
rect 11057 10044 11069 10047
rect 9732 10016 11069 10044
rect 9732 10004 9738 10016
rect 11057 10013 11069 10016
rect 11103 10044 11115 10047
rect 11146 10044 11152 10056
rect 11103 10016 11152 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12452 10016 12909 10044
rect 2133 9979 2191 9985
rect 2133 9945 2145 9979
rect 2179 9976 2191 9979
rect 2866 9976 2872 9988
rect 2179 9948 2872 9976
rect 2179 9945 2191 9948
rect 2133 9939 2191 9945
rect 2866 9936 2872 9948
rect 2924 9936 2930 9988
rect 4884 9979 4942 9985
rect 4884 9945 4896 9979
rect 4930 9976 4942 9979
rect 5258 9976 5264 9988
rect 4930 9948 5264 9976
rect 4930 9945 4942 9948
rect 4884 9939 4942 9945
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 6822 9985 6828 9988
rect 6816 9976 6828 9985
rect 6783 9948 6828 9976
rect 6816 9939 6828 9948
rect 6822 9936 6828 9939
rect 6880 9936 6886 9988
rect 8570 9936 8576 9988
rect 8628 9976 8634 9988
rect 11330 9985 11336 9988
rect 9370 9979 9428 9985
rect 9370 9976 9382 9979
rect 8628 9948 9382 9976
rect 8628 9936 8634 9948
rect 9370 9945 9382 9948
rect 9416 9945 9428 9979
rect 9370 9939 9428 9945
rect 11324 9939 11336 9985
rect 11330 9936 11336 9939
rect 11388 9936 11394 9988
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6730 9908 6736 9920
rect 6052 9880 6736 9908
rect 6052 9868 6058 9880
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12452 9917 12480 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 12989 9979 13047 9985
rect 12989 9976 13001 9979
rect 12584 9948 13001 9976
rect 12584 9936 12590 9948
rect 12989 9945 13001 9948
rect 13035 9945 13047 9979
rect 12989 9939 13047 9945
rect 13170 9936 13176 9988
rect 13228 9936 13234 9988
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 13780 9948 14289 9976
rect 13780 9936 13786 9948
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 14476 9976 14504 10075
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 16577 10115 16635 10121
rect 16577 10112 16589 10115
rect 15304 10084 16589 10112
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10044 14611 10047
rect 14918 10044 14924 10056
rect 14599 10016 14924 10044
rect 14599 10013 14611 10016
rect 14553 10007 14611 10013
rect 14918 10004 14924 10016
rect 14976 10044 14982 10056
rect 15304 10053 15332 10084
rect 16577 10081 16589 10084
rect 16623 10112 16635 10115
rect 17494 10112 17500 10124
rect 16623 10084 17500 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 20898 10072 20904 10124
rect 20956 10072 20962 10124
rect 23382 10072 23388 10124
rect 23440 10072 23446 10124
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 14976 10016 15301 10044
rect 14976 10004 14982 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15562 10044 15568 10056
rect 15289 10007 15347 10013
rect 15397 10016 15568 10044
rect 15102 9976 15108 9988
rect 14476 9948 15108 9976
rect 14277 9939 14335 9945
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 12437 9911 12495 9917
rect 12437 9908 12449 9911
rect 11940 9880 12449 9908
rect 11940 9868 11946 9880
rect 12437 9877 12449 9880
rect 12483 9877 12495 9911
rect 12437 9871 12495 9877
rect 12894 9868 12900 9920
rect 12952 9868 12958 9920
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15397 9908 15425 10016
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 16482 10004 16488 10056
rect 16540 10004 16546 10056
rect 16776 10016 17724 10044
rect 15068 9880 15425 9908
rect 15473 9911 15531 9917
rect 15068 9868 15074 9880
rect 15473 9877 15485 9911
rect 15519 9908 15531 9911
rect 16776 9908 16804 10016
rect 17696 9985 17724 10016
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 18380 10016 19625 10044
rect 18380 10004 18386 10016
rect 19613 10013 19625 10016
rect 19659 10044 19671 10047
rect 20346 10044 20352 10056
rect 19659 10016 20352 10044
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 23400 10044 23428 10072
rect 22603 10016 23428 10044
rect 23845 10047 23903 10053
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 23952 10044 23980 10152
rect 26786 10140 26792 10152
rect 26844 10140 26850 10192
rect 27982 10140 27988 10192
rect 28040 10180 28046 10192
rect 28040 10152 28580 10180
rect 28040 10140 28046 10152
rect 25501 10115 25559 10121
rect 25501 10081 25513 10115
rect 25547 10112 25559 10115
rect 27157 10115 27215 10121
rect 27157 10112 27169 10115
rect 25547 10084 27169 10112
rect 25547 10081 25559 10084
rect 25501 10075 25559 10081
rect 27157 10081 27169 10084
rect 27203 10081 27215 10115
rect 27157 10075 27215 10081
rect 27798 10072 27804 10124
rect 27856 10112 27862 10124
rect 28552 10121 28580 10152
rect 28445 10115 28503 10121
rect 28445 10112 28457 10115
rect 27856 10084 28457 10112
rect 27856 10072 27862 10084
rect 28445 10081 28457 10084
rect 28491 10081 28503 10115
rect 28445 10075 28503 10081
rect 28537 10115 28595 10121
rect 28537 10081 28549 10115
rect 28583 10081 28595 10115
rect 28537 10075 28595 10081
rect 29454 10072 29460 10124
rect 29512 10112 29518 10124
rect 30006 10112 30012 10124
rect 29512 10084 30012 10112
rect 29512 10072 29518 10084
rect 30006 10072 30012 10084
rect 30064 10112 30070 10124
rect 30193 10115 30251 10121
rect 30193 10112 30205 10115
rect 30064 10084 30205 10112
rect 30064 10072 30070 10084
rect 30193 10081 30205 10084
rect 30239 10081 30251 10115
rect 30193 10075 30251 10081
rect 30926 10072 30932 10124
rect 30984 10072 30990 10124
rect 31772 10112 31800 10208
rect 31312 10084 31800 10112
rect 23891 10016 23980 10044
rect 24029 10047 24087 10053
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 17681 9979 17739 9985
rect 16868 9948 17632 9976
rect 16868 9917 16896 9948
rect 15519 9880 16804 9908
rect 16853 9911 16911 9917
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 16853 9877 16865 9911
rect 16899 9877 16911 9911
rect 16853 9871 16911 9877
rect 17310 9868 17316 9920
rect 17368 9868 17374 9920
rect 17494 9917 17500 9920
rect 17481 9911 17500 9917
rect 17481 9877 17493 9911
rect 17481 9871 17500 9877
rect 17494 9868 17500 9871
rect 17552 9868 17558 9920
rect 17604 9908 17632 9948
rect 17681 9945 17693 9979
rect 17727 9976 17739 9979
rect 18230 9976 18236 9988
rect 17727 9948 18236 9976
rect 17727 9945 17739 9948
rect 17681 9939 17739 9945
rect 18230 9936 18236 9948
rect 18288 9976 18294 9988
rect 18877 9979 18935 9985
rect 18877 9976 18889 9979
rect 18288 9948 18889 9976
rect 18288 9936 18294 9948
rect 18877 9945 18889 9948
rect 18923 9945 18935 9979
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 18877 9939 18935 9945
rect 19536 9948 19717 9976
rect 18667 9911 18725 9917
rect 18667 9908 18679 9911
rect 17604 9880 18679 9908
rect 18667 9877 18679 9880
rect 18713 9908 18725 9911
rect 19242 9908 19248 9920
rect 18713 9880 19248 9908
rect 18713 9877 18725 9880
rect 18667 9871 18725 9877
rect 19242 9868 19248 9880
rect 19300 9908 19306 9920
rect 19536 9908 19564 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 19705 9939 19763 9945
rect 23198 9936 23204 9988
rect 23256 9936 23262 9988
rect 23385 9979 23443 9985
rect 23385 9945 23397 9979
rect 23431 9976 23443 9979
rect 23658 9976 23664 9988
rect 23431 9948 23664 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 23658 9936 23664 9948
rect 23716 9976 23722 9988
rect 24044 9976 24072 10007
rect 24946 10004 24952 10056
rect 25004 10053 25010 10056
rect 25004 10047 25040 10053
rect 25028 10013 25040 10047
rect 25004 10007 25040 10013
rect 25004 10004 25010 10007
rect 25406 10004 25412 10056
rect 25464 10004 25470 10056
rect 26050 10004 26056 10056
rect 26108 10044 26114 10056
rect 26145 10047 26203 10053
rect 26145 10044 26157 10047
rect 26108 10016 26157 10044
rect 26108 10004 26114 10016
rect 26145 10013 26157 10016
rect 26191 10013 26203 10047
rect 26145 10007 26203 10013
rect 26326 10004 26332 10056
rect 26384 10004 26390 10056
rect 26510 10004 26516 10056
rect 26568 10004 26574 10056
rect 27341 10047 27399 10053
rect 27341 10013 27353 10047
rect 27387 10013 27399 10047
rect 27341 10007 27399 10013
rect 23716 9948 24072 9976
rect 26237 9979 26295 9985
rect 23716 9936 23722 9948
rect 26237 9945 26249 9979
rect 26283 9976 26295 9979
rect 26602 9976 26608 9988
rect 26283 9948 26608 9976
rect 26283 9945 26295 9948
rect 26237 9939 26295 9945
rect 26602 9936 26608 9948
rect 26660 9936 26666 9988
rect 27356 9976 27384 10007
rect 27430 10004 27436 10056
rect 27488 10004 27494 10056
rect 27706 10004 27712 10056
rect 27764 10004 27770 10056
rect 28258 10004 28264 10056
rect 28316 10044 28322 10056
rect 28353 10047 28411 10053
rect 28353 10044 28365 10047
rect 28316 10016 28365 10044
rect 28316 10004 28322 10016
rect 28353 10013 28365 10016
rect 28399 10013 28411 10047
rect 28353 10007 28411 10013
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10044 28687 10047
rect 28718 10044 28724 10056
rect 28675 10016 28724 10044
rect 28675 10013 28687 10016
rect 28629 10007 28687 10013
rect 28718 10004 28724 10016
rect 28776 10044 28782 10056
rect 30098 10044 30104 10056
rect 28776 10016 30104 10044
rect 28776 10004 28782 10016
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 31110 10004 31116 10056
rect 31168 10004 31174 10056
rect 31312 10053 31340 10084
rect 31297 10047 31355 10053
rect 31297 10013 31309 10047
rect 31343 10013 31355 10047
rect 31297 10007 31355 10013
rect 31757 10047 31815 10053
rect 31757 10013 31769 10047
rect 31803 10013 31815 10047
rect 31757 10007 31815 10013
rect 27356 9948 28212 9976
rect 19300 9880 19564 9908
rect 19300 9868 19306 9880
rect 19794 9868 19800 9920
rect 19852 9868 19858 9920
rect 24854 9868 24860 9920
rect 24912 9868 24918 9920
rect 25038 9868 25044 9920
rect 25096 9868 25102 9920
rect 25958 9868 25964 9920
rect 26016 9868 26022 9920
rect 27614 9868 27620 9920
rect 27672 9908 27678 9920
rect 27982 9908 27988 9920
rect 27672 9880 27988 9908
rect 27672 9868 27678 9880
rect 27982 9868 27988 9880
rect 28040 9868 28046 9920
rect 28184 9917 28212 9948
rect 30834 9936 30840 9988
rect 30892 9936 30898 9988
rect 31772 9976 31800 10007
rect 31938 10004 31944 10056
rect 31996 10004 32002 10056
rect 31036 9948 31800 9976
rect 28169 9911 28227 9917
rect 28169 9877 28181 9911
rect 28215 9908 28227 9911
rect 29733 9911 29791 9917
rect 29733 9908 29745 9911
rect 28215 9880 29745 9908
rect 28215 9877 28227 9880
rect 28169 9871 28227 9877
rect 29733 9877 29745 9880
rect 29779 9877 29791 9911
rect 29733 9871 29791 9877
rect 30377 9911 30435 9917
rect 30377 9877 30389 9911
rect 30423 9908 30435 9911
rect 31036 9908 31064 9948
rect 30423 9880 31064 9908
rect 30423 9877 30435 9880
rect 30377 9871 30435 9877
rect 1104 9818 32632 9840
rect 1104 9766 8792 9818
rect 8844 9766 8856 9818
rect 8908 9766 8920 9818
rect 8972 9766 8984 9818
rect 9036 9766 9048 9818
rect 9100 9766 16634 9818
rect 16686 9766 16698 9818
rect 16750 9766 16762 9818
rect 16814 9766 16826 9818
rect 16878 9766 16890 9818
rect 16942 9766 24476 9818
rect 24528 9766 24540 9818
rect 24592 9766 24604 9818
rect 24656 9766 24668 9818
rect 24720 9766 24732 9818
rect 24784 9766 32318 9818
rect 32370 9766 32382 9818
rect 32434 9766 32446 9818
rect 32498 9766 32510 9818
rect 32562 9766 32574 9818
rect 32626 9766 32632 9818
rect 1104 9744 32632 9766
rect 1949 9707 2007 9713
rect 1949 9673 1961 9707
rect 1995 9704 2007 9707
rect 2314 9704 2320 9716
rect 1995 9676 2320 9704
rect 1995 9673 2007 9676
rect 1949 9667 2007 9673
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2409 9707 2467 9713
rect 2409 9673 2421 9707
rect 2455 9673 2467 9707
rect 6086 9704 6092 9716
rect 2409 9667 2467 9673
rect 4448 9676 6092 9704
rect 1581 9639 1639 9645
rect 1581 9605 1593 9639
rect 1627 9605 1639 9639
rect 1581 9599 1639 9605
rect 1797 9639 1855 9645
rect 1797 9605 1809 9639
rect 1843 9636 1855 9639
rect 2424 9636 2452 9667
rect 1843 9608 2452 9636
rect 1843 9605 1855 9608
rect 1797 9599 1855 9605
rect 1596 9568 1624 9599
rect 2222 9568 2228 9580
rect 1596 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2424 9500 2452 9608
rect 3421 9639 3479 9645
rect 3421 9605 3433 9639
rect 3467 9636 3479 9639
rect 4341 9639 4399 9645
rect 4341 9636 4353 9639
rect 3467 9608 4353 9636
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 4341 9605 4353 9608
rect 4387 9605 4399 9639
rect 4341 9599 4399 9605
rect 2774 9528 2780 9580
rect 2832 9528 2838 9580
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3108 9540 3648 9568
rect 3108 9528 3114 9540
rect 2685 9503 2743 9509
rect 2424 9472 2636 9500
rect 2608 9432 2636 9472
rect 2685 9469 2697 9503
rect 2731 9500 2743 9503
rect 3068 9500 3096 9528
rect 2731 9472 3096 9500
rect 3421 9503 3479 9509
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 3421 9469 3433 9503
rect 3467 9469 3479 9503
rect 3620 9500 3648 9540
rect 3694 9528 3700 9580
rect 3752 9528 3758 9580
rect 4154 9528 4160 9580
rect 4212 9528 4218 9580
rect 4448 9577 4476 9676
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 14369 9707 14427 9713
rect 6604 9676 6960 9704
rect 6604 9664 6610 9676
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 4540 9608 6009 9636
rect 4540 9577 4568 9608
rect 5997 9605 6009 9608
rect 6043 9636 6055 9639
rect 6362 9636 6368 9648
rect 6043 9608 6368 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 6932 9580 6960 9676
rect 14369 9673 14381 9707
rect 14415 9704 14427 9707
rect 14550 9704 14556 9716
rect 14415 9676 14556 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 18524 9676 19472 9704
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 9525 9639 9583 9645
rect 9364 9608 9444 9636
rect 9364 9596 9370 9608
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 4448 9500 4476 9531
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7173 9571 7231 9577
rect 7173 9568 7185 9571
rect 7064 9540 7185 9568
rect 7064 9528 7070 9540
rect 7173 9537 7185 9540
rect 7219 9537 7231 9571
rect 9416 9568 9444 9608
rect 9525 9605 9537 9639
rect 9571 9636 9583 9639
rect 12894 9636 12900 9648
rect 9571 9608 12900 9636
rect 9571 9605 9583 9608
rect 9525 9599 9583 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 14458 9636 14464 9648
rect 13004 9608 14464 9636
rect 9674 9568 9680 9580
rect 9416 9540 9680 9568
rect 7173 9531 7231 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9568 10563 9571
rect 11882 9568 11888 9580
rect 10551 9540 11888 9568
rect 10551 9537 10563 9540
rect 10505 9531 10563 9537
rect 3620 9472 4476 9500
rect 5629 9503 5687 9509
rect 3421 9463 3479 9469
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 5902 9500 5908 9512
rect 5675 9472 5908 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 3050 9432 3056 9444
rect 2608 9404 3056 9432
rect 3050 9392 3056 9404
rect 3108 9432 3114 9444
rect 3436 9432 3464 9463
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10520 9500 10548 9531
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12618 9568 12624 9580
rect 12207 9540 12624 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 10008 9472 10548 9500
rect 10781 9503 10839 9509
rect 10008 9460 10014 9472
rect 10781 9469 10793 9503
rect 10827 9500 10839 9503
rect 11330 9500 11336 9512
rect 10827 9472 11336 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 12084 9500 12112 9531
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13004 9577 13032 9608
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 15194 9596 15200 9648
rect 15252 9596 15258 9648
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9636 16359 9639
rect 17126 9636 17132 9648
rect 16347 9608 17132 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 18524 9636 18552 9676
rect 17460 9608 18552 9636
rect 18601 9639 18659 9645
rect 17460 9596 17466 9608
rect 18601 9605 18613 9639
rect 18647 9636 18659 9639
rect 19334 9636 19340 9648
rect 18647 9608 19340 9636
rect 18647 9605 18659 9608
rect 18601 9599 18659 9605
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 19444 9636 19472 9676
rect 19794 9664 19800 9716
rect 19852 9704 19858 9716
rect 20441 9707 20499 9713
rect 20441 9704 20453 9707
rect 19852 9676 20453 9704
rect 19852 9664 19858 9676
rect 20441 9673 20453 9676
rect 20487 9673 20499 9707
rect 20441 9667 20499 9673
rect 22186 9664 22192 9716
rect 22244 9664 22250 9716
rect 25038 9664 25044 9716
rect 25096 9704 25102 9716
rect 25409 9707 25467 9713
rect 25409 9704 25421 9707
rect 25096 9676 25421 9704
rect 25096 9664 25102 9676
rect 25409 9673 25421 9676
rect 25455 9704 25467 9707
rect 26050 9704 26056 9716
rect 25455 9676 26056 9704
rect 25455 9673 25467 9676
rect 25409 9667 25467 9673
rect 26050 9664 26056 9676
rect 26108 9664 26114 9716
rect 26344 9676 27844 9704
rect 19610 9636 19616 9648
rect 19444 9608 19616 9636
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 21910 9636 21916 9648
rect 20824 9608 21916 9636
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9568 13047 9571
rect 13078 9568 13084 9580
rect 13035 9540 13084 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13262 9577 13268 9580
rect 13256 9568 13268 9577
rect 13223 9540 13268 9568
rect 13256 9531 13268 9540
rect 13262 9528 13268 9531
rect 13320 9528 13326 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14660 9540 15025 9568
rect 12526 9500 12532 9512
rect 12084 9472 12532 9500
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 11701 9435 11759 9441
rect 11701 9432 11713 9435
rect 3108 9404 3464 9432
rect 9508 9404 11713 9432
rect 3108 9392 3114 9404
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 2958 9364 2964 9376
rect 1811 9336 2964 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 3605 9367 3663 9373
rect 3605 9364 3617 9367
rect 3200 9336 3617 9364
rect 3200 9324 3206 9336
rect 3605 9333 3617 9336
rect 3651 9333 3663 9367
rect 3605 9327 3663 9333
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 9508 9373 9536 9404
rect 11701 9401 11713 9404
rect 11747 9401 11759 9435
rect 11701 9395 11759 9401
rect 14660 9432 14688 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9568 15347 9571
rect 15470 9568 15476 9580
rect 15335 9540 15476 9568
rect 15335 9537 15347 9540
rect 15289 9531 15347 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 17310 9568 17316 9580
rect 16163 9540 17316 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 18230 9528 18236 9580
rect 18288 9568 18294 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 18288 9540 18337 9568
rect 18288 9528 18294 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 19242 9528 19248 9580
rect 19300 9528 19306 9580
rect 19426 9528 19432 9580
rect 19484 9528 19490 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 20824 9577 20852 9608
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22554 9636 22560 9648
rect 22204 9608 22560 9636
rect 22204 9577 22232 9608
rect 22554 9596 22560 9608
rect 22612 9636 22618 9648
rect 23658 9636 23664 9648
rect 22612 9608 23664 9636
rect 22612 9596 22618 9608
rect 23658 9596 23664 9608
rect 23716 9596 23722 9648
rect 25314 9596 25320 9648
rect 25372 9636 25378 9648
rect 26142 9636 26148 9648
rect 25372 9608 26148 9636
rect 25372 9596 25378 9608
rect 26142 9596 26148 9608
rect 26200 9596 26206 9648
rect 26234 9596 26240 9648
rect 26292 9636 26298 9648
rect 26344 9636 26372 9676
rect 26292 9608 26372 9636
rect 26453 9639 26511 9645
rect 26292 9596 26298 9608
rect 26453 9605 26465 9639
rect 26499 9636 26511 9639
rect 26602 9636 26608 9648
rect 26499 9608 26608 9636
rect 26499 9605 26511 9608
rect 26453 9599 26511 9605
rect 26602 9596 26608 9608
rect 26660 9596 26666 9648
rect 26694 9596 26700 9648
rect 26752 9636 26758 9648
rect 27246 9636 27252 9648
rect 26752 9608 27252 9636
rect 26752 9596 26758 9608
rect 27246 9596 27252 9608
rect 27304 9636 27310 9648
rect 27304 9608 27752 9636
rect 27304 9596 27310 9608
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9537 20867 9571
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 20809 9531 20867 9537
rect 20916 9540 22017 9568
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15378 9500 15384 9512
rect 15252 9472 15384 9500
rect 15252 9460 15258 9472
rect 15378 9460 15384 9472
rect 15436 9500 15442 9512
rect 15930 9500 15936 9512
rect 15436 9472 15936 9500
rect 15436 9460 15442 9472
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 18601 9503 18659 9509
rect 18601 9469 18613 9503
rect 18647 9500 18659 9503
rect 19061 9503 19119 9509
rect 19061 9500 19073 9503
rect 18647 9472 19073 9500
rect 18647 9469 18659 9472
rect 18601 9463 18659 9469
rect 19061 9469 19073 9472
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 20438 9500 20444 9512
rect 19392 9472 20444 9500
rect 19392 9460 19398 9472
rect 20438 9460 20444 9472
rect 20496 9500 20502 9512
rect 20717 9503 20775 9509
rect 20717 9500 20729 9503
rect 20496 9472 20729 9500
rect 20496 9460 20502 9472
rect 20717 9469 20729 9472
rect 20763 9469 20775 9503
rect 20717 9463 20775 9469
rect 17310 9432 17316 9444
rect 14660 9404 17316 9432
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 7616 9336 8309 9364
rect 7616 9324 7622 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 8297 9327 8355 9333
rect 9493 9367 9551 9373
rect 9493 9333 9505 9367
rect 9539 9333 9551 9367
rect 9493 9327 9551 9333
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 11606 9364 11612 9376
rect 9723 9336 11612 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 14660 9364 14688 9404
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 18380 9404 18429 9432
rect 18380 9392 18386 9404
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 20916 9432 20944 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 22916 9571 22974 9577
rect 22916 9537 22928 9571
rect 22962 9568 22974 9571
rect 24302 9568 24308 9580
rect 22962 9540 24308 9568
rect 22962 9537 22974 9540
rect 22916 9531 22974 9537
rect 24302 9528 24308 9540
rect 24360 9528 24366 9580
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 24964 9540 27537 9568
rect 24964 9512 24992 9540
rect 27525 9537 27537 9540
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 27614 9528 27620 9580
rect 27672 9528 27678 9580
rect 22649 9503 22707 9509
rect 22649 9500 22661 9503
rect 22066 9472 22661 9500
rect 18417 9395 18475 9401
rect 19352 9404 20944 9432
rect 12032 9336 14688 9364
rect 12032 9324 12038 9336
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14792 9336 14841 9364
rect 14792 9324 14798 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 19352 9364 19380 9404
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 21910 9432 21916 9444
rect 21140 9404 21916 9432
rect 21140 9392 21146 9404
rect 21910 9392 21916 9404
rect 21968 9432 21974 9444
rect 22066 9432 22094 9472
rect 22649 9469 22661 9472
rect 22695 9469 22707 9503
rect 24946 9500 24952 9512
rect 22649 9463 22707 9469
rect 24044 9472 24952 9500
rect 24044 9441 24072 9472
rect 24946 9460 24952 9472
rect 25004 9460 25010 9512
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 27632 9500 27660 9528
rect 25639 9472 27660 9500
rect 27724 9500 27752 9608
rect 27816 9568 27844 9676
rect 27890 9664 27896 9716
rect 27948 9704 27954 9716
rect 29454 9704 29460 9716
rect 27948 9676 29460 9704
rect 27948 9664 27954 9676
rect 29454 9664 29460 9676
rect 29512 9664 29518 9716
rect 30466 9664 30472 9716
rect 30524 9664 30530 9716
rect 31110 9664 31116 9716
rect 31168 9704 31174 9716
rect 31665 9707 31723 9713
rect 31665 9704 31677 9707
rect 31168 9676 31677 9704
rect 31168 9664 31174 9676
rect 31665 9673 31677 9676
rect 31711 9673 31723 9707
rect 31665 9667 31723 9673
rect 28905 9639 28963 9645
rect 28905 9636 28917 9639
rect 28460 9608 28917 9636
rect 28166 9568 28172 9580
rect 27816 9540 28172 9568
rect 28166 9528 28172 9540
rect 28224 9528 28230 9580
rect 28460 9500 28488 9608
rect 28905 9605 28917 9608
rect 28951 9636 28963 9639
rect 30484 9636 30512 9664
rect 28951 9608 30512 9636
rect 30552 9639 30610 9645
rect 28951 9605 28963 9608
rect 28905 9599 28963 9605
rect 30552 9605 30564 9639
rect 30598 9636 30610 9639
rect 30834 9636 30840 9648
rect 30598 9608 30840 9636
rect 30598 9605 30610 9608
rect 30552 9599 30610 9605
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 28537 9571 28595 9577
rect 28537 9537 28549 9571
rect 28583 9537 28595 9571
rect 28537 9531 28595 9537
rect 28721 9571 28779 9577
rect 28721 9537 28733 9571
rect 28767 9537 28779 9571
rect 28721 9531 28779 9537
rect 27724 9472 28488 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 21968 9404 22094 9432
rect 24029 9435 24087 9441
rect 21968 9392 21974 9404
rect 24029 9401 24041 9435
rect 24075 9401 24087 9435
rect 24029 9395 24087 9401
rect 24688 9404 25084 9432
rect 17184 9336 19380 9364
rect 17184 9324 17190 9336
rect 19610 9324 19616 9376
rect 19668 9364 19674 9376
rect 24688 9364 24716 9404
rect 19668 9336 24716 9364
rect 19668 9324 19674 9336
rect 24762 9324 24768 9376
rect 24820 9364 24826 9376
rect 24949 9367 25007 9373
rect 24949 9364 24961 9367
rect 24820 9336 24961 9364
rect 24820 9324 24826 9336
rect 24949 9333 24961 9336
rect 24995 9333 25007 9367
rect 25056 9364 25084 9404
rect 26142 9392 26148 9444
rect 26200 9432 26206 9444
rect 28552 9432 28580 9531
rect 26200 9404 28580 9432
rect 28736 9432 28764 9531
rect 28810 9528 28816 9580
rect 28868 9568 28874 9580
rect 29365 9571 29423 9577
rect 29365 9568 29377 9571
rect 28868 9540 29377 9568
rect 28868 9528 28874 9540
rect 29365 9537 29377 9540
rect 29411 9537 29423 9571
rect 29365 9531 29423 9537
rect 29454 9528 29460 9580
rect 29512 9528 29518 9580
rect 30282 9528 30288 9580
rect 30340 9528 30346 9580
rect 29641 9503 29699 9509
rect 29641 9469 29653 9503
rect 29687 9500 29699 9503
rect 29730 9500 29736 9512
rect 29687 9472 29736 9500
rect 29687 9469 29699 9472
rect 29641 9463 29699 9469
rect 29730 9460 29736 9472
rect 29788 9460 29794 9512
rect 28736 9404 29868 9432
rect 26200 9392 26206 9404
rect 26234 9364 26240 9376
rect 25056 9336 26240 9364
rect 24949 9327 25007 9333
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 26421 9367 26479 9373
rect 26421 9333 26433 9367
rect 26467 9364 26479 9367
rect 26510 9364 26516 9376
rect 26467 9336 26516 9364
rect 26467 9333 26479 9336
rect 26421 9327 26479 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 26605 9367 26663 9373
rect 26605 9333 26617 9367
rect 26651 9364 26663 9367
rect 26786 9364 26792 9376
rect 26651 9336 26792 9364
rect 26651 9333 26663 9336
rect 26605 9327 26663 9333
rect 26786 9324 26792 9336
rect 26844 9324 26850 9376
rect 27709 9367 27767 9373
rect 27709 9333 27721 9367
rect 27755 9364 27767 9367
rect 27798 9364 27804 9376
rect 27755 9336 27804 9364
rect 27755 9333 27767 9336
rect 27709 9327 27767 9333
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 27890 9324 27896 9376
rect 27948 9364 27954 9376
rect 28736 9364 28764 9404
rect 27948 9336 28764 9364
rect 29549 9367 29607 9373
rect 27948 9324 27954 9336
rect 29549 9333 29561 9367
rect 29595 9364 29607 9367
rect 29730 9364 29736 9376
rect 29595 9336 29736 9364
rect 29595 9333 29607 9336
rect 29549 9327 29607 9333
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 29840 9364 29868 9404
rect 31478 9364 31484 9376
rect 29840 9336 31484 9364
rect 31478 9324 31484 9336
rect 31536 9324 31542 9376
rect 1104 9274 32476 9296
rect 1104 9222 4871 9274
rect 4923 9222 4935 9274
rect 4987 9222 4999 9274
rect 5051 9222 5063 9274
rect 5115 9222 5127 9274
rect 5179 9222 12713 9274
rect 12765 9222 12777 9274
rect 12829 9222 12841 9274
rect 12893 9222 12905 9274
rect 12957 9222 12969 9274
rect 13021 9222 20555 9274
rect 20607 9222 20619 9274
rect 20671 9222 20683 9274
rect 20735 9222 20747 9274
rect 20799 9222 20811 9274
rect 20863 9222 28397 9274
rect 28449 9222 28461 9274
rect 28513 9222 28525 9274
rect 28577 9222 28589 9274
rect 28641 9222 28653 9274
rect 28705 9222 32476 9274
rect 1104 9200 32476 9222
rect 3421 9163 3479 9169
rect 3421 9129 3433 9163
rect 3467 9160 3479 9163
rect 4154 9160 4160 9172
rect 3467 9132 4160 9160
rect 3467 9129 3479 9132
rect 3421 9123 3479 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 5718 9120 5724 9172
rect 5776 9160 5782 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5776 9132 5825 9160
rect 5776 9120 5782 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 6512 9132 6561 9160
rect 6512 9120 6518 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 10226 9160 10232 9172
rect 10091 9132 10232 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12676 9132 13001 9160
rect 12676 9120 12682 9132
rect 12989 9129 13001 9132
rect 13035 9160 13047 9163
rect 13170 9160 13176 9172
rect 13035 9132 13176 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 16022 9160 16028 9172
rect 13740 9132 16028 9160
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 3142 9092 3148 9104
rect 2455 9064 3148 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 3234 9052 3240 9104
rect 3292 9052 3298 9104
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 7558 9092 7564 9104
rect 3568 9064 7564 9092
rect 3568 9052 3574 9064
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 1995 8996 2912 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2038 8916 2044 8968
rect 2096 8916 2102 8968
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2774 8956 2780 8968
rect 2280 8928 2780 8956
rect 2280 8916 2286 8928
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 2884 8888 2912 8996
rect 3050 8984 3056 9036
rect 3108 8984 3114 9036
rect 3252 9024 3280 9052
rect 3160 8996 3280 9024
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3160 8956 3188 8996
rect 3007 8928 3188 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3694 8956 3700 8968
rect 3292 8928 3700 8956
rect 3292 8916 3298 8928
rect 3694 8916 3700 8928
rect 3752 8956 3758 8968
rect 4172 8965 4200 9064
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9092 8539 9095
rect 9122 9092 9128 9104
rect 8527 9064 9128 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 9916 9064 10701 9092
rect 9916 9052 9922 9064
rect 10689 9061 10701 9064
rect 10735 9092 10747 9095
rect 10870 9092 10876 9104
rect 10735 9064 10876 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 10870 9052 10876 9064
rect 10928 9052 10934 9104
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 13740 9092 13768 9132
rect 16022 9120 16028 9132
rect 16080 9160 16086 9172
rect 16080 9132 17724 9160
rect 16080 9120 16086 9132
rect 13688 9064 13768 9092
rect 13688 9052 13694 9064
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7282 9024 7288 9036
rect 6963 8996 7288 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 13078 9024 13084 9036
rect 7392 8996 9444 9024
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3752 8928 3985 8956
rect 3752 8916 3758 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 2884 8860 3004 8888
rect 2976 8832 3004 8860
rect 3326 8848 3332 8900
rect 3384 8888 3390 8900
rect 4264 8888 4292 8919
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 7392 8965 7420 8996
rect 9416 8968 9444 8996
rect 12084 8996 13084 9024
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 4764 8928 6745 8956
rect 4764 8916 4770 8928
rect 6733 8925 6745 8928
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7377 8919 7435 8925
rect 7484 8928 7757 8956
rect 4614 8888 4620 8900
rect 3384 8860 4620 8888
rect 3384 8848 3390 8860
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5442 8848 5448 8900
rect 5500 8848 5506 8900
rect 5626 8848 5632 8900
rect 5684 8848 5690 8900
rect 6638 8848 6644 8900
rect 6696 8888 6702 8900
rect 7484 8888 7512 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 6696 8860 7512 8888
rect 7561 8891 7619 8897
rect 6696 8848 6702 8860
rect 7561 8857 7573 8891
rect 7607 8857 7619 8891
rect 7561 8851 7619 8857
rect 2958 8780 2964 8832
rect 3016 8780 3022 8832
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 7576 8820 7604 8851
rect 7650 8848 7656 8900
rect 7708 8848 7714 8900
rect 7760 8888 7788 8919
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 8352 8928 8401 8956
rect 8352 8916 8358 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8536 8928 8585 8956
rect 8536 8916 8542 8928
rect 8573 8925 8585 8928
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9456 8928 9505 8956
rect 9456 8916 9462 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9493 8919 9551 8925
rect 9600 8928 9873 8956
rect 9600 8888 9628 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 7760 8860 9628 8888
rect 9674 8848 9680 8900
rect 9732 8848 9738 8900
rect 9769 8891 9827 8897
rect 9769 8857 9781 8891
rect 9815 8857 9827 8891
rect 9876 8888 9904 8919
rect 11790 8916 11796 8968
rect 11848 8965 11854 8968
rect 11848 8956 11860 8965
rect 11848 8928 11893 8956
rect 11848 8919 11860 8928
rect 11848 8916 11854 8919
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 12084 8965 12112 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 12032 8928 12081 8956
rect 12032 8916 12038 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12710 8956 12716 8968
rect 12492 8928 12716 8956
rect 12492 8916 12498 8928
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12768 8928 12817 8956
rect 12768 8916 12774 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 13740 8965 13768 9064
rect 15841 9095 15899 9101
rect 15841 9061 15853 9095
rect 15887 9092 15899 9095
rect 17586 9092 17592 9104
rect 15887 9064 17592 9092
rect 15887 9061 15899 9064
rect 15841 9055 15899 9061
rect 17586 9052 17592 9064
rect 17644 9052 17650 9104
rect 17696 9092 17724 9132
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18288 9132 18705 9160
rect 18288 9120 18294 9132
rect 18693 9129 18705 9132
rect 18739 9160 18751 9163
rect 19334 9160 19340 9172
rect 18739 9132 19340 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 20809 9163 20867 9169
rect 20809 9160 20821 9163
rect 19484 9132 20821 9160
rect 19484 9120 19490 9132
rect 20809 9129 20821 9132
rect 20855 9129 20867 9163
rect 20809 9123 20867 9129
rect 18506 9092 18512 9104
rect 17696 9064 18512 9092
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 14458 8984 14464 9036
rect 14516 8984 14522 9036
rect 20824 9024 20852 9123
rect 26602 9120 26608 9172
rect 26660 9120 26666 9172
rect 27065 9163 27123 9169
rect 27065 9160 27077 9163
rect 26712 9132 27077 9160
rect 26142 9052 26148 9104
rect 26200 9092 26206 9104
rect 26712 9092 26740 9132
rect 27065 9129 27077 9132
rect 27111 9129 27123 9163
rect 27065 9123 27123 9129
rect 28994 9120 29000 9172
rect 29052 9160 29058 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 29052 9132 29837 9160
rect 29052 9120 29058 9132
rect 29825 9129 29837 9132
rect 29871 9129 29883 9163
rect 29825 9123 29883 9129
rect 27617 9095 27675 9101
rect 27617 9092 27629 9095
rect 26200 9064 26740 9092
rect 26804 9064 27629 9092
rect 26200 9052 26206 9064
rect 16316 8996 19380 9024
rect 20824 8996 21496 9024
rect 14734 8965 14740 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13504 8928 13553 8956
rect 13504 8916 13510 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 14728 8956 14740 8965
rect 14695 8928 14740 8956
rect 13725 8919 13783 8925
rect 14728 8919 14740 8928
rect 14734 8916 14740 8919
rect 14792 8916 14798 8968
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 16316 8965 16344 8996
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 15160 8928 16313 8956
rect 15160 8916 15166 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 17034 8956 17040 8968
rect 16531 8928 17040 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 12158 8888 12164 8900
rect 9876 8860 12164 8888
rect 9769 8851 9827 8857
rect 3108 8792 7604 8820
rect 3108 8780 3114 8792
rect 7926 8780 7932 8832
rect 7984 8780 7990 8832
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 9784 8820 9812 8851
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 12621 8891 12679 8897
rect 12621 8888 12633 8891
rect 12400 8860 12633 8888
rect 12400 8848 12406 8860
rect 12621 8857 12633 8860
rect 12667 8857 12679 8891
rect 12621 8851 12679 8857
rect 13633 8891 13691 8897
rect 13633 8857 13645 8891
rect 13679 8888 13691 8891
rect 17126 8888 17132 8900
rect 13679 8860 17132 8888
rect 13679 8857 13691 8860
rect 13633 8851 13691 8857
rect 10042 8820 10048 8832
rect 8168 8792 10048 8820
rect 8168 8780 8174 8792
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 13648 8820 13676 8851
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 18506 8848 18512 8900
rect 18564 8848 18570 8900
rect 19352 8888 19380 8996
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 20898 8956 20904 8968
rect 19475 8928 20904 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 21468 8965 21496 8996
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 23532 8996 24593 9024
rect 23532 8984 23538 8996
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24581 8987 24639 8993
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 19696 8891 19754 8897
rect 19352 8860 19656 8888
rect 19628 8832 19656 8860
rect 19696 8857 19708 8891
rect 19742 8888 19754 8891
rect 19886 8888 19892 8900
rect 19742 8860 19892 8888
rect 19742 8857 19754 8860
rect 19696 8851 19754 8857
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 20438 8848 20444 8900
rect 20496 8888 20502 8900
rect 21284 8888 21312 8919
rect 21910 8916 21916 8968
rect 21968 8956 21974 8968
rect 22462 8965 22468 8968
rect 22189 8959 22247 8965
rect 22189 8956 22201 8959
rect 21968 8928 22201 8956
rect 21968 8916 21974 8928
rect 22189 8925 22201 8928
rect 22235 8925 22247 8959
rect 22456 8956 22468 8965
rect 22423 8928 22468 8956
rect 22189 8919 22247 8925
rect 22456 8919 22468 8928
rect 22462 8916 22468 8919
rect 22520 8916 22526 8968
rect 24762 8916 24768 8968
rect 24820 8916 24826 8968
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 20496 8860 21312 8888
rect 20496 8848 20502 8860
rect 21358 8848 21364 8900
rect 21416 8888 21422 8900
rect 25884 8888 25912 8919
rect 25958 8916 25964 8968
rect 26016 8916 26022 8968
rect 26234 8956 26240 8968
rect 26068 8928 26240 8956
rect 26068 8888 26096 8928
rect 26234 8916 26240 8928
rect 26292 8916 26298 8968
rect 26804 8965 26832 9064
rect 27617 9061 27629 9064
rect 27663 9061 27675 9095
rect 28905 9095 28963 9101
rect 28905 9092 28917 9095
rect 27617 9055 27675 9061
rect 28092 9064 28917 9092
rect 27706 8984 27712 9036
rect 27764 9024 27770 9036
rect 28092 9033 28120 9064
rect 28905 9061 28917 9064
rect 28951 9061 28963 9095
rect 28905 9055 28963 9061
rect 28077 9027 28135 9033
rect 28077 9024 28089 9027
rect 27764 8996 28089 9024
rect 27764 8984 27770 8996
rect 28077 8993 28089 8996
rect 28123 8993 28135 9027
rect 28077 8987 28135 8993
rect 28166 8984 28172 9036
rect 28224 8984 28230 9036
rect 29638 8984 29644 9036
rect 29696 9024 29702 9036
rect 29696 8996 29960 9024
rect 29696 8984 29702 8996
rect 26789 8959 26847 8965
rect 26789 8925 26801 8959
rect 26835 8925 26847 8959
rect 26789 8919 26847 8925
rect 26881 8959 26939 8965
rect 26881 8925 26893 8959
rect 26927 8956 26939 8959
rect 26970 8956 26976 8968
rect 26927 8928 26976 8956
rect 26927 8925 26939 8928
rect 26881 8919 26939 8925
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 27798 8956 27804 8968
rect 27203 8928 27804 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8956 28043 8959
rect 28718 8956 28724 8968
rect 28031 8928 28724 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 28718 8916 28724 8928
rect 28776 8956 28782 8968
rect 28813 8959 28871 8965
rect 28813 8956 28825 8959
rect 28776 8928 28825 8956
rect 28776 8916 28782 8928
rect 28813 8925 28825 8928
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 28902 8916 28908 8968
rect 28960 8956 28966 8968
rect 28997 8959 29055 8965
rect 28997 8956 29009 8959
rect 28960 8928 29009 8956
rect 28960 8916 28966 8928
rect 28997 8925 29009 8928
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29730 8916 29736 8968
rect 29788 8916 29794 8968
rect 29932 8965 29960 8996
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8925 29975 8959
rect 29917 8919 29975 8925
rect 30561 8959 30619 8965
rect 30561 8925 30573 8959
rect 30607 8925 30619 8959
rect 30561 8919 30619 8925
rect 21416 8860 25820 8888
rect 25884 8860 26096 8888
rect 26145 8891 26203 8897
rect 21416 8848 21422 8860
rect 25792 8832 25820 8860
rect 26145 8857 26157 8891
rect 26191 8888 26203 8891
rect 30576 8888 30604 8919
rect 26191 8860 30604 8888
rect 26191 8857 26203 8860
rect 26145 8851 26203 8857
rect 10284 8792 13676 8820
rect 10284 8780 10290 8792
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 16264 8792 16313 8820
rect 16264 8780 16270 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 18690 8820 18696 8832
rect 18748 8829 18754 8832
rect 18748 8823 18767 8829
rect 17276 8792 18696 8820
rect 17276 8780 17282 8792
rect 18690 8780 18696 8792
rect 18755 8789 18767 8823
rect 18748 8783 18767 8789
rect 18877 8823 18935 8829
rect 18877 8789 18889 8823
rect 18923 8820 18935 8823
rect 19426 8820 19432 8832
rect 18923 8792 19432 8820
rect 18923 8789 18935 8792
rect 18877 8783 18935 8789
rect 18748 8780 18754 8783
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 19610 8780 19616 8832
rect 19668 8820 19674 8832
rect 22002 8820 22008 8832
rect 19668 8792 22008 8820
rect 19668 8780 19674 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 23569 8823 23627 8829
rect 23569 8789 23581 8823
rect 23615 8820 23627 8823
rect 23658 8820 23664 8832
rect 23615 8792 23664 8820
rect 23615 8789 23627 8792
rect 23569 8783 23627 8789
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 24949 8823 25007 8829
rect 24949 8789 24961 8823
rect 24995 8820 25007 8823
rect 25222 8820 25228 8832
rect 24995 8792 25228 8820
rect 24995 8789 25007 8792
rect 24949 8783 25007 8789
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 25774 8780 25780 8832
rect 25832 8820 25838 8832
rect 27890 8820 27896 8832
rect 25832 8792 27896 8820
rect 25832 8780 25838 8792
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 30374 8780 30380 8832
rect 30432 8780 30438 8832
rect 1104 8730 32632 8752
rect 1104 8678 8792 8730
rect 8844 8678 8856 8730
rect 8908 8678 8920 8730
rect 8972 8678 8984 8730
rect 9036 8678 9048 8730
rect 9100 8678 16634 8730
rect 16686 8678 16698 8730
rect 16750 8678 16762 8730
rect 16814 8678 16826 8730
rect 16878 8678 16890 8730
rect 16942 8678 24476 8730
rect 24528 8678 24540 8730
rect 24592 8678 24604 8730
rect 24656 8678 24668 8730
rect 24720 8678 24732 8730
rect 24784 8678 32318 8730
rect 32370 8678 32382 8730
rect 32434 8678 32446 8730
rect 32498 8678 32510 8730
rect 32562 8678 32574 8730
rect 32626 8678 32632 8730
rect 1104 8656 32632 8678
rect 2961 8619 3019 8625
rect 2961 8585 2973 8619
rect 3007 8616 3019 8619
rect 3050 8616 3056 8628
rect 3007 8588 3056 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 5736 8588 7757 8616
rect 3421 8551 3479 8557
rect 3421 8548 3433 8551
rect 2056 8520 3433 8548
rect 2056 8492 2084 8520
rect 3421 8517 3433 8520
rect 3467 8517 3479 8551
rect 3421 8511 3479 8517
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 5736 8548 5764 8588
rect 7745 8585 7757 8588
rect 7791 8616 7803 8619
rect 8386 8616 8392 8628
rect 7791 8588 8392 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 9861 8619 9919 8625
rect 8680 8588 9720 8616
rect 4672 8520 5764 8548
rect 4672 8508 4678 8520
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 8478 8548 8484 8560
rect 7340 8520 8484 8548
rect 7340 8508 7346 8520
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2038 8480 2044 8492
rect 1995 8452 2044 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 1780 8344 1808 8443
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 2774 8480 2780 8492
rect 2639 8452 2780 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 3384 8452 3617 8480
rect 3384 8440 3390 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 5718 8440 5724 8492
rect 5776 8440 5782 8492
rect 5994 8480 6000 8492
rect 5828 8452 6000 8480
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 1903 8384 2513 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 5534 8412 5540 8424
rect 3936 8384 5540 8412
rect 3936 8372 3942 8384
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 2958 8344 2964 8356
rect 1780 8316 2964 8344
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 5828 8344 5856 8452
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6420 8452 6561 8480
rect 6420 8440 6426 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7708 8452 7849 8480
rect 7708 8440 7714 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 7984 8452 8585 8480
rect 7984 8440 7990 8452
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8412 5963 8415
rect 8680 8412 8708 8588
rect 9692 8548 9720 8588
rect 9861 8585 9873 8619
rect 9907 8616 9919 8619
rect 10318 8616 10324 8628
rect 9907 8588 10324 8616
rect 9907 8585 9919 8588
rect 9861 8579 9919 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10965 8619 11023 8625
rect 10965 8585 10977 8619
rect 11011 8616 11023 8619
rect 12526 8616 12532 8628
rect 11011 8588 12532 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 12526 8576 12532 8588
rect 12584 8616 12590 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 12584 8588 12633 8616
rect 12584 8576 12590 8588
rect 12621 8585 12633 8588
rect 12667 8585 12679 8619
rect 12621 8579 12679 8585
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 14642 8616 14648 8628
rect 13504 8588 14648 8616
rect 13504 8576 13510 8588
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 14918 8576 14924 8628
rect 14976 8576 14982 8628
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 19889 8619 19947 8625
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 20254 8616 20260 8628
rect 19935 8588 20260 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 22370 8576 22376 8628
rect 22428 8576 22434 8628
rect 24302 8576 24308 8628
rect 24360 8576 24366 8628
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 26513 8619 26571 8625
rect 24452 8588 25176 8616
rect 24452 8576 24458 8588
rect 10226 8548 10232 8560
rect 9692 8520 10232 8548
rect 9692 8489 9720 8520
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 10928 8520 11560 8548
rect 10928 8508 10934 8520
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 9950 8480 9956 8492
rect 9907 8452 9956 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8480 10563 8483
rect 11532 8480 11560 8520
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11664 8520 11713 8548
rect 11664 8508 11670 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 12342 8548 12348 8560
rect 11701 8511 11759 8517
rect 11900 8520 12348 8548
rect 11900 8489 11928 8520
rect 12342 8508 12348 8520
rect 12400 8548 12406 8560
rect 12400 8520 12572 8548
rect 12400 8508 12406 8520
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 10551 8452 11468 8480
rect 11532 8452 11897 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 5951 8384 8708 8412
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9766 8412 9772 8424
rect 8812 8384 9772 8412
rect 8812 8372 8818 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9968 8412 9996 8440
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 9968 8384 10609 8412
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 11440 8412 11468 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12158 8480 12164 8492
rect 12023 8452 12164 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12544 8489 12572 8520
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 14516 8520 16344 8548
rect 14516 8508 14522 8520
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12710 8440 12716 8492
rect 12768 8440 12774 8492
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13311 8452 13921 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 15102 8480 15108 8492
rect 14240 8452 15108 8480
rect 14240 8440 14246 8452
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 16045 8483 16103 8489
rect 16045 8449 16057 8483
rect 16091 8480 16103 8483
rect 16206 8480 16212 8492
rect 16091 8452 16212 8480
rect 16091 8449 16103 8452
rect 16045 8443 16103 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16316 8489 16344 8520
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 21358 8548 21364 8560
rect 18564 8520 21364 8548
rect 18564 8508 18570 8520
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 24412 8548 24440 8576
rect 23768 8520 24440 8548
rect 25148 8548 25176 8588
rect 26513 8585 26525 8619
rect 26559 8616 26571 8619
rect 27614 8616 27620 8628
rect 26559 8588 27620 8616
rect 26559 8585 26571 8588
rect 26513 8579 26571 8585
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 29822 8576 29828 8628
rect 29880 8616 29886 8628
rect 30929 8619 30987 8625
rect 30929 8616 30941 8619
rect 29880 8588 30941 8616
rect 29880 8576 29886 8588
rect 30929 8585 30941 8588
rect 30975 8585 30987 8619
rect 30929 8579 30987 8585
rect 30282 8548 30288 8560
rect 25148 8520 30288 8548
rect 17494 8489 17500 8492
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16347 8452 17233 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17488 8443 17500 8489
rect 17494 8440 17500 8443
rect 17552 8440 17558 8492
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 20714 8480 20720 8492
rect 18748 8452 20720 8480
rect 18748 8440 18754 8452
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 21013 8483 21071 8489
rect 21013 8449 21025 8483
rect 21059 8480 21071 8483
rect 21174 8480 21180 8492
rect 21059 8452 21180 8480
rect 21059 8449 21071 8452
rect 21013 8443 21071 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21910 8480 21916 8492
rect 21315 8452 21916 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21910 8440 21916 8452
rect 21968 8440 21974 8492
rect 23474 8440 23480 8492
rect 23532 8489 23538 8492
rect 23768 8489 23796 8520
rect 23532 8443 23544 8489
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24854 8480 24860 8492
rect 24443 8452 24860 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 23532 8440 23538 8443
rect 12618 8412 12624 8424
rect 11440 8384 12624 8412
rect 10597 8375 10655 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 3844 8316 5856 8344
rect 5920 8316 7052 8344
rect 3844 8304 3850 8316
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 5920 8276 5948 8316
rect 5776 8248 5948 8276
rect 5776 8236 5782 8248
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 6733 8279 6791 8285
rect 6733 8276 6745 8279
rect 6696 8248 6745 8276
rect 6696 8236 6702 8248
rect 6733 8245 6745 8248
rect 6779 8245 6791 8279
rect 7024 8276 7052 8316
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 8389 8347 8447 8353
rect 8389 8344 8401 8347
rect 7156 8316 8401 8344
rect 7156 8304 7162 8316
rect 8389 8313 8401 8316
rect 8435 8313 8447 8347
rect 11606 8344 11612 8356
rect 8389 8307 8447 8313
rect 8496 8316 11612 8344
rect 8496 8276 8524 8316
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 11698 8304 11704 8356
rect 11756 8304 11762 8356
rect 13449 8347 13507 8353
rect 13449 8313 13461 8347
rect 13495 8344 13507 8347
rect 14550 8344 14556 8356
rect 13495 8316 14556 8344
rect 13495 8313 13507 8316
rect 13449 8307 13507 8313
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 7024 8248 8524 8276
rect 6733 8239 6791 8245
rect 10318 8236 10324 8288
rect 10376 8276 10382 8288
rect 10962 8276 10968 8288
rect 10376 8248 10968 8276
rect 10376 8236 10382 8248
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 17218 8276 17224 8288
rect 14700 8248 17224 8276
rect 14700 8236 14706 8248
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 24228 8276 24256 8443
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 25148 8489 25176 8520
rect 25406 8489 25412 8492
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 25400 8443 25412 8489
rect 25406 8440 25412 8443
rect 25464 8440 25470 8492
rect 27172 8489 27200 8520
rect 27157 8483 27215 8489
rect 27157 8449 27169 8483
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27246 8440 27252 8492
rect 27304 8480 27310 8492
rect 29564 8489 29592 8520
rect 30282 8508 30288 8520
rect 30340 8508 30346 8560
rect 27413 8483 27471 8489
rect 27413 8480 27425 8483
rect 27304 8452 27425 8480
rect 27304 8440 27310 8452
rect 27413 8449 27425 8452
rect 27459 8449 27471 8483
rect 27413 8443 27471 8449
rect 29549 8483 29607 8489
rect 29549 8449 29561 8483
rect 29595 8449 29607 8483
rect 29549 8443 29607 8449
rect 29816 8483 29874 8489
rect 29816 8449 29828 8483
rect 29862 8480 29874 8483
rect 30374 8480 30380 8492
rect 29862 8452 30380 8480
rect 29862 8449 29874 8452
rect 29816 8443 29874 8449
rect 30374 8440 30380 8452
rect 30432 8440 30438 8492
rect 24762 8276 24768 8288
rect 23624 8248 24768 8276
rect 23624 8236 23630 8248
rect 24762 8236 24768 8248
rect 24820 8236 24826 8288
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 28537 8279 28595 8285
rect 28537 8276 28549 8279
rect 27856 8248 28549 8276
rect 27856 8236 27862 8248
rect 28537 8245 28549 8248
rect 28583 8245 28595 8279
rect 28537 8239 28595 8245
rect 1104 8186 32476 8208
rect 1104 8134 4871 8186
rect 4923 8134 4935 8186
rect 4987 8134 4999 8186
rect 5051 8134 5063 8186
rect 5115 8134 5127 8186
rect 5179 8134 12713 8186
rect 12765 8134 12777 8186
rect 12829 8134 12841 8186
rect 12893 8134 12905 8186
rect 12957 8134 12969 8186
rect 13021 8134 20555 8186
rect 20607 8134 20619 8186
rect 20671 8134 20683 8186
rect 20735 8134 20747 8186
rect 20799 8134 20811 8186
rect 20863 8134 28397 8186
rect 28449 8134 28461 8186
rect 28513 8134 28525 8186
rect 28577 8134 28589 8186
rect 28641 8134 28653 8186
rect 28705 8134 32476 8186
rect 1104 8112 32476 8134
rect 2774 8032 2780 8084
rect 2832 8032 2838 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 7006 8072 7012 8084
rect 6779 8044 7012 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8352 8044 8585 8072
rect 8352 8032 8358 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 9490 8072 9496 8084
rect 9355 8044 9496 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17034 8072 17040 8084
rect 16991 8044 17040 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 17552 8044 17601 8072
rect 17552 8032 17558 8044
rect 17589 8041 17601 8044
rect 17635 8041 17647 8075
rect 17589 8035 17647 8041
rect 19886 8032 19892 8084
rect 19944 8032 19950 8084
rect 20640 8044 21128 8072
rect 10226 7964 10232 8016
rect 10284 7964 10290 8016
rect 17402 7964 17408 8016
rect 17460 7964 17466 8016
rect 20640 8004 20668 8044
rect 17512 7976 20668 8004
rect 20717 8007 20775 8013
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7936 5963 7939
rect 6914 7936 6920 7948
rect 5951 7908 6920 7936
rect 5951 7905 5963 7908
rect 5905 7899 5963 7905
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6972 7908 7205 7936
rect 6972 7896 6978 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 14458 7896 14464 7948
rect 14516 7896 14522 7948
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 17034 7936 17040 7948
rect 16807 7908 17040 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 17034 7896 17040 7908
rect 17092 7936 17098 7948
rect 17420 7936 17448 7964
rect 17092 7908 17448 7936
rect 17092 7896 17098 7908
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2866 7868 2872 7880
rect 2823 7840 2872 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3234 7868 3240 7880
rect 3007 7840 3240 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7098 7868 7104 7880
rect 6595 7840 7104 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 9950 7868 9956 7880
rect 9416 7840 9956 7868
rect 5660 7803 5718 7809
rect 5660 7769 5672 7803
rect 5706 7800 5718 7803
rect 6362 7800 6368 7812
rect 5706 7772 6368 7800
rect 5706 7769 5718 7772
rect 5660 7763 5718 7769
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7438 7803 7496 7809
rect 7438 7800 7450 7803
rect 7064 7772 7450 7800
rect 7064 7760 7070 7772
rect 7438 7769 7450 7772
rect 7484 7769 7496 7803
rect 7438 7763 7496 7769
rect 9293 7803 9351 7809
rect 9293 7769 9305 7803
rect 9339 7800 9351 7803
rect 9416 7800 9444 7840
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 11112 7840 11161 7868
rect 11112 7828 11118 7840
rect 11149 7837 11161 7840
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 11882 7868 11888 7880
rect 11839 7840 11888 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 14717 7871 14775 7877
rect 14717 7868 14729 7871
rect 14608 7840 14729 7868
rect 14608 7828 14614 7840
rect 14717 7837 14729 7840
rect 14763 7837 14775 7871
rect 14717 7831 14775 7837
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 17126 7868 17132 7880
rect 16715 7840 17132 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 17368 7840 17417 7868
rect 17368 7828 17374 7840
rect 17405 7837 17417 7840
rect 17451 7868 17463 7871
rect 17512 7868 17540 7976
rect 20717 7973 20729 8007
rect 20763 7973 20775 8007
rect 20717 7967 20775 7973
rect 19426 7896 19432 7948
rect 19484 7896 19490 7948
rect 17451 7840 17540 7868
rect 17589 7871 17647 7877
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17862 7868 17868 7880
rect 17635 7840 17868 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19668 7840 19717 7868
rect 19668 7828 19674 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 20732 7868 20760 7967
rect 21100 7936 21128 8044
rect 21174 8032 21180 8084
rect 21232 8032 21238 8084
rect 23566 8072 23572 8084
rect 22066 8044 23572 8072
rect 22066 7936 22094 8044
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 23661 8075 23719 8081
rect 23661 8041 23673 8075
rect 23707 8072 23719 8075
rect 24302 8072 24308 8084
rect 23707 8044 24308 8072
rect 23707 8041 23719 8044
rect 23661 8035 23719 8041
rect 24302 8032 24308 8044
rect 24360 8032 24366 8084
rect 25406 8032 25412 8084
rect 25464 8032 25470 8084
rect 26973 8075 27031 8081
rect 26973 8041 26985 8075
rect 27019 8072 27031 8075
rect 27246 8072 27252 8084
rect 27019 8044 27252 8072
rect 27019 8041 27031 8044
rect 26973 8035 27031 8041
rect 27246 8032 27252 8044
rect 27304 8032 27310 8084
rect 27985 8075 28043 8081
rect 27985 8041 27997 8075
rect 28031 8072 28043 8075
rect 28166 8072 28172 8084
rect 28031 8044 28172 8072
rect 28031 8041 28043 8044
rect 27985 8035 28043 8041
rect 28166 8032 28172 8044
rect 28224 8032 28230 8084
rect 23017 8007 23075 8013
rect 23017 7973 23029 8007
rect 23063 7973 23075 8007
rect 23017 7967 23075 7973
rect 21100 7908 22094 7936
rect 21376 7877 21404 7908
rect 22370 7896 22376 7948
rect 22428 7936 22434 7948
rect 22554 7936 22560 7948
rect 22428 7908 22560 7936
rect 22428 7896 22434 7908
rect 22554 7896 22560 7908
rect 22612 7936 22618 7948
rect 22612 7908 22876 7936
rect 22612 7896 22618 7908
rect 22848 7877 22876 7908
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20732 7840 21189 7868
rect 20441 7831 20499 7837
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 21361 7871 21419 7877
rect 21361 7837 21373 7871
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 23032 7868 23060 7967
rect 23474 7964 23480 8016
rect 23532 8004 23538 8016
rect 24581 8007 24639 8013
rect 24581 8004 24593 8007
rect 23532 7976 24593 8004
rect 23532 7964 23538 7976
rect 24581 7973 24593 7976
rect 24627 7973 24639 8007
rect 24581 7967 24639 7973
rect 27709 7939 27767 7945
rect 27709 7905 27721 7939
rect 27755 7936 27767 7939
rect 27798 7936 27804 7948
rect 27755 7908 27804 7936
rect 27755 7905 27767 7908
rect 27709 7899 27767 7905
rect 27798 7896 27804 7908
rect 27856 7896 27862 7948
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23032 7840 24593 7868
rect 22833 7831 22891 7837
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 9339 7772 9444 7800
rect 9493 7803 9551 7809
rect 9339 7769 9351 7772
rect 9293 7763 9351 7769
rect 9493 7769 9505 7803
rect 9539 7769 9551 7803
rect 9493 7763 9551 7769
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3878 7732 3884 7744
rect 2924 7704 3884 7732
rect 2924 7692 2930 7704
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4525 7735 4583 7741
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 5258 7732 5264 7744
rect 4571 7704 5264 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 7190 7732 7196 7744
rect 6788 7704 7196 7732
rect 6788 7692 6794 7704
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8720 7704 9137 7732
rect 8720 7692 8726 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9125 7695 9183 7701
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 9508 7732 9536 7763
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 10229 7803 10287 7809
rect 10229 7800 10241 7803
rect 10192 7772 10241 7800
rect 10192 7760 10198 7772
rect 10229 7769 10241 7772
rect 10275 7769 10287 7803
rect 10229 7763 10287 7769
rect 11241 7803 11299 7809
rect 11241 7769 11253 7803
rect 11287 7800 11299 7803
rect 12038 7803 12096 7809
rect 12038 7800 12050 7803
rect 11287 7772 12050 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 12038 7769 12050 7772
rect 12084 7769 12096 7803
rect 12038 7763 12096 7769
rect 15378 7760 15384 7812
rect 15436 7800 15442 7812
rect 16301 7803 16359 7809
rect 16301 7800 16313 7803
rect 15436 7772 16313 7800
rect 15436 7760 15442 7772
rect 16301 7769 16313 7772
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 16390 7760 16396 7812
rect 16448 7760 16454 7812
rect 17678 7760 17684 7812
rect 17736 7800 17742 7812
rect 20456 7800 20484 7831
rect 20717 7803 20775 7809
rect 17736 7772 20668 7800
rect 17736 7760 17742 7772
rect 9456 7704 9536 7732
rect 9456 7692 9462 7704
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 9640 7704 10057 7732
rect 9640 7692 9646 7704
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 13170 7692 13176 7744
rect 13228 7732 13234 7744
rect 13722 7732 13728 7744
rect 13228 7704 13728 7732
rect 13228 7692 13234 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 13872 7704 15853 7732
rect 13872 7692 13878 7704
rect 15841 7701 15853 7704
rect 15887 7732 15899 7735
rect 15930 7732 15936 7744
rect 15887 7704 15936 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 20254 7692 20260 7744
rect 20312 7732 20318 7744
rect 20533 7735 20591 7741
rect 20533 7732 20545 7735
rect 20312 7704 20545 7732
rect 20312 7692 20318 7704
rect 20533 7701 20545 7704
rect 20579 7701 20591 7735
rect 20640 7732 20668 7772
rect 20717 7769 20729 7803
rect 20763 7800 20775 7803
rect 22370 7800 22376 7812
rect 20763 7772 22376 7800
rect 20763 7769 20775 7772
rect 20717 7763 20775 7769
rect 22370 7760 22376 7772
rect 22428 7760 22434 7812
rect 22756 7732 22784 7831
rect 24762 7828 24768 7880
rect 24820 7828 24826 7880
rect 25222 7828 25228 7880
rect 25280 7828 25286 7880
rect 26786 7828 26792 7880
rect 26844 7828 26850 7880
rect 27614 7828 27620 7880
rect 27672 7828 27678 7880
rect 23017 7803 23075 7809
rect 23017 7769 23029 7803
rect 23063 7769 23075 7803
rect 23017 7763 23075 7769
rect 20640 7704 22784 7732
rect 23032 7732 23060 7763
rect 23290 7760 23296 7812
rect 23348 7800 23354 7812
rect 23845 7803 23903 7809
rect 23845 7800 23857 7803
rect 23348 7772 23857 7800
rect 23348 7760 23354 7772
rect 23845 7769 23857 7772
rect 23891 7769 23903 7803
rect 23845 7763 23903 7769
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 23032 7704 23489 7732
rect 20533 7695 20591 7701
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 23645 7735 23703 7741
rect 23645 7701 23657 7735
rect 23691 7732 23703 7735
rect 24394 7732 24400 7744
rect 23691 7704 24400 7732
rect 23691 7701 23703 7704
rect 23645 7695 23703 7701
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 1104 7642 32632 7664
rect 1104 7590 8792 7642
rect 8844 7590 8856 7642
rect 8908 7590 8920 7642
rect 8972 7590 8984 7642
rect 9036 7590 9048 7642
rect 9100 7590 16634 7642
rect 16686 7590 16698 7642
rect 16750 7590 16762 7642
rect 16814 7590 16826 7642
rect 16878 7590 16890 7642
rect 16942 7590 24476 7642
rect 24528 7590 24540 7642
rect 24592 7590 24604 7642
rect 24656 7590 24668 7642
rect 24720 7590 24732 7642
rect 24784 7590 32318 7642
rect 32370 7590 32382 7642
rect 32434 7590 32446 7642
rect 32498 7590 32510 7642
rect 32562 7590 32574 7642
rect 32626 7590 32632 7642
rect 1104 7568 32632 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 2958 7528 2964 7540
rect 2915 7500 2964 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 4433 7531 4491 7537
rect 3108 7500 4108 7528
rect 3108 7488 3114 7500
rect 2240 7432 3004 7460
rect 2240 7401 2268 7432
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2866 7392 2872 7404
rect 2455 7364 2872 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 2976 7324 3004 7432
rect 4080 7401 4108 7500
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 5626 7528 5632 7540
rect 4479 7500 5632 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 7006 7528 7012 7540
rect 6871 7500 7012 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 5828 7460 5856 7491
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9490 7488 9496 7540
rect 9548 7488 9554 7540
rect 9968 7500 10824 7528
rect 6638 7460 6644 7472
rect 5828 7432 6644 7460
rect 6638 7420 6644 7432
rect 6696 7460 6702 7472
rect 7653 7463 7711 7469
rect 6696 7432 7420 7460
rect 6696 7420 6702 7432
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5718 7392 5724 7404
rect 5491 7364 5724 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5816 7395 5874 7401
rect 5816 7361 5828 7395
rect 5862 7361 5874 7395
rect 5816 7355 5874 7361
rect 3234 7324 3240 7336
rect 2976 7296 3240 7324
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 4154 7284 4160 7336
rect 4212 7284 4218 7336
rect 5350 7284 5356 7336
rect 5408 7284 5414 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5828 7324 5856 7355
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 7392 7401 7420 7432
rect 7653 7429 7665 7463
rect 7699 7460 7711 7463
rect 8662 7460 8668 7472
rect 7699 7432 8668 7460
rect 7699 7429 7711 7432
rect 7653 7423 7711 7429
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 9140 7460 9168 7488
rect 9398 7460 9404 7472
rect 9140 7432 9404 7460
rect 9398 7420 9404 7432
rect 9456 7460 9462 7472
rect 9582 7460 9588 7472
rect 9456 7432 9588 7460
rect 9456 7420 9462 7432
rect 9582 7420 9588 7432
rect 9640 7460 9646 7472
rect 9968 7469 9996 7500
rect 9953 7463 10011 7469
rect 9953 7460 9965 7463
rect 9640 7432 9965 7460
rect 9640 7420 9646 7432
rect 9953 7429 9965 7432
rect 9999 7429 10011 7463
rect 9953 7423 10011 7429
rect 10134 7420 10140 7472
rect 10192 7469 10198 7472
rect 10192 7463 10211 7469
rect 10199 7429 10211 7463
rect 10192 7423 10211 7429
rect 10192 7420 10198 7423
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7392 7527 7395
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7515 7364 8125 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 8113 7361 8125 7364
rect 8159 7392 8171 7395
rect 8294 7392 8300 7404
rect 8159 7364 8300 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 5592 7296 5856 7324
rect 6932 7324 6960 7355
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9766 7392 9772 7404
rect 9355 7364 9772 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9048 7324 9076 7355
rect 9766 7352 9772 7364
rect 9824 7392 9830 7404
rect 10318 7392 10324 7404
rect 9824 7364 10324 7392
rect 9824 7352 9830 7364
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10796 7401 10824 7500
rect 11330 7488 11336 7540
rect 11388 7528 11394 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11388 7500 12173 7528
rect 11388 7488 11394 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 12308 7500 12357 7528
rect 12308 7488 12314 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 11020 7432 11069 7460
rect 11020 7420 11026 7432
rect 11057 7429 11069 7432
rect 11103 7429 11115 7463
rect 12360 7460 12388 7491
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16390 7528 16396 7540
rect 16347 7500 16396 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 17862 7488 17868 7540
rect 17920 7488 17926 7540
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19576 7500 19993 7528
rect 19576 7488 19582 7500
rect 19981 7497 19993 7500
rect 20027 7497 20039 7531
rect 19981 7491 20039 7497
rect 20149 7531 20207 7537
rect 20149 7497 20161 7531
rect 20195 7528 20207 7531
rect 21634 7528 21640 7540
rect 20195 7500 21640 7528
rect 20195 7497 20207 7500
rect 20149 7491 20207 7497
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 22741 7531 22799 7537
rect 22741 7497 22753 7531
rect 22787 7528 22799 7531
rect 23845 7531 23903 7537
rect 23845 7528 23857 7531
rect 22787 7500 23857 7528
rect 22787 7497 22799 7500
rect 22741 7491 22799 7497
rect 23845 7497 23857 7500
rect 23891 7497 23903 7531
rect 23845 7491 23903 7497
rect 17696 7460 17724 7488
rect 12360 7432 17724 7460
rect 20349 7463 20407 7469
rect 11057 7423 11115 7429
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7361 10931 7395
rect 12250 7392 12256 7404
rect 12308 7401 12314 7404
rect 12308 7395 12344 7401
rect 12244 7364 12256 7392
rect 10873 7355 10931 7361
rect 9582 7324 9588 7336
rect 6932 7296 7696 7324
rect 9048 7296 9588 7324
rect 5592 7284 5598 7296
rect 3326 7256 3332 7268
rect 2746 7228 3332 7256
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2746 7188 2774 7228
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 3421 7259 3479 7265
rect 3421 7225 3433 7259
rect 3467 7256 3479 7259
rect 4246 7256 4252 7268
rect 3467 7228 4252 7256
rect 3467 7225 3479 7228
rect 3421 7219 3479 7225
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 7668 7265 7696 7296
rect 9582 7284 9588 7296
rect 9640 7324 9646 7336
rect 10888 7324 10916 7355
rect 12250 7352 12256 7364
rect 12332 7392 12344 7395
rect 13170 7392 13176 7404
rect 12332 7364 13176 7392
rect 12332 7361 12344 7364
rect 12308 7355 12344 7361
rect 12308 7352 12314 7355
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 13722 7352 13728 7404
rect 13780 7352 13786 7404
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 13924 7401 13952 7432
rect 20349 7429 20361 7463
rect 20395 7460 20407 7463
rect 22646 7460 22652 7472
rect 20395 7432 22652 7460
rect 20395 7429 20407 7432
rect 20349 7423 20407 7429
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 16117 7395 16175 7401
rect 15427 7364 15884 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 9640 7296 10916 7324
rect 9640 7284 9646 7296
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 11664 7296 12725 7324
rect 11664 7284 11670 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13078 7324 13084 7336
rect 12851 7296 13084 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 7653 7259 7711 7265
rect 7653 7225 7665 7259
rect 7699 7225 7711 7259
rect 7653 7219 7711 7225
rect 8110 7216 8116 7268
rect 8168 7256 8174 7268
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 8168 7228 8217 7256
rect 8168 7216 8174 7228
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 8205 7219 8263 7225
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 10781 7259 10839 7265
rect 10781 7256 10793 7259
rect 10008 7228 10793 7256
rect 10008 7216 10014 7228
rect 2363 7160 2774 7188
rect 3053 7191 3111 7197
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 4430 7188 4436 7200
rect 3099 7160 4436 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 5997 7191 6055 7197
rect 5997 7157 6009 7191
rect 6043 7188 6055 7191
rect 6546 7188 6552 7200
rect 6043 7160 6552 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 8570 7148 8576 7200
rect 8628 7148 8634 7200
rect 10152 7197 10180 7228
rect 10781 7225 10793 7228
rect 10827 7225 10839 7259
rect 12728 7256 12756 7287
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 13446 7256 13452 7268
rect 12728 7228 13452 7256
rect 10781 7219 10839 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 15212 7256 15240 7355
rect 15856 7333 15884 7364
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 17740 7395 17798 7401
rect 16163 7364 17632 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 15887 7296 16436 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 16408 7256 16436 7296
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 17310 7284 17316 7336
rect 17368 7284 17374 7336
rect 17604 7324 17632 7364
rect 17740 7361 17752 7395
rect 17786 7392 17798 7395
rect 18598 7392 18604 7404
rect 17786 7364 18604 7392
rect 17786 7361 17798 7364
rect 17740 7355 17798 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 20364 7324 20392 7423
rect 22646 7420 22652 7432
rect 22704 7420 22710 7472
rect 23860 7460 23888 7491
rect 24302 7488 24308 7540
rect 24360 7488 24366 7540
rect 24394 7488 24400 7540
rect 24452 7528 24458 7540
rect 25225 7531 25283 7537
rect 25225 7528 25237 7531
rect 24452 7500 25237 7528
rect 24452 7488 24458 7500
rect 25225 7497 25237 7500
rect 25271 7497 25283 7531
rect 25225 7491 25283 7497
rect 24673 7463 24731 7469
rect 24673 7460 24685 7463
rect 23860 7432 24685 7460
rect 24673 7429 24685 7432
rect 24719 7460 24731 7463
rect 25317 7463 25375 7469
rect 25317 7460 25329 7463
rect 24719 7432 25329 7460
rect 24719 7429 24731 7432
rect 24673 7423 24731 7429
rect 25317 7429 25329 7432
rect 25363 7429 25375 7463
rect 25317 7423 25375 7429
rect 22554 7352 22560 7404
rect 22612 7352 22618 7404
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7392 23443 7395
rect 24489 7395 24547 7401
rect 23431 7364 24440 7392
rect 23431 7361 23443 7364
rect 23385 7355 23443 7361
rect 17604 7296 20392 7324
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 20496 7296 20821 7324
rect 20496 7284 20502 7296
rect 20809 7293 20821 7296
rect 20855 7324 20867 7327
rect 22756 7324 22784 7355
rect 23014 7324 23020 7336
rect 20855 7296 23020 7324
rect 20855 7293 20867 7296
rect 20809 7287 20867 7293
rect 23014 7284 23020 7296
rect 23072 7284 23078 7336
rect 23477 7327 23535 7333
rect 23477 7293 23489 7327
rect 23523 7293 23535 7327
rect 24412 7324 24440 7364
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24578 7392 24584 7404
rect 24535 7364 24584 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24578 7352 24584 7364
rect 24636 7352 24642 7404
rect 24765 7395 24823 7401
rect 24765 7392 24777 7395
rect 24688 7364 24777 7392
rect 24688 7324 24716 7364
rect 24765 7361 24777 7364
rect 24811 7361 24823 7395
rect 24765 7355 24823 7361
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 25225 7395 25283 7401
rect 25225 7392 25237 7395
rect 24912 7364 25237 7392
rect 24912 7352 24918 7364
rect 25225 7361 25237 7364
rect 25271 7361 25283 7395
rect 25225 7355 25283 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 24412 7296 24716 7324
rect 23477 7287 23535 7293
rect 17954 7256 17960 7268
rect 15212 7228 15976 7256
rect 16408 7228 17960 7256
rect 10137 7191 10195 7197
rect 10137 7157 10149 7191
rect 10183 7157 10195 7191
rect 10137 7151 10195 7157
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 10410 7188 10416 7200
rect 10367 7160 10416 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 15948 7197 15976 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 21085 7259 21143 7265
rect 21085 7256 21097 7259
rect 20312 7228 21097 7256
rect 20312 7216 20318 7228
rect 21085 7225 21097 7228
rect 21131 7256 21143 7259
rect 22462 7256 22468 7268
rect 21131 7228 22468 7256
rect 21131 7225 21143 7228
rect 21085 7219 21143 7225
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 23201 7259 23259 7265
rect 23201 7256 23213 7259
rect 22572 7228 23213 7256
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 17126 7188 17132 7200
rect 15979 7160 17132 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 20165 7191 20223 7197
rect 20165 7157 20177 7191
rect 20211 7188 20223 7191
rect 20438 7188 20444 7200
rect 20211 7160 20444 7188
rect 20211 7157 20223 7160
rect 20165 7151 20223 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 21269 7191 21327 7197
rect 21269 7188 21281 7191
rect 21232 7160 21281 7188
rect 21232 7148 21238 7160
rect 21269 7157 21281 7160
rect 21315 7157 21327 7191
rect 21269 7151 21327 7157
rect 21726 7148 21732 7200
rect 21784 7188 21790 7200
rect 22572 7188 22600 7228
rect 23201 7225 23213 7228
rect 23247 7225 23259 7259
rect 23492 7256 23520 7287
rect 24688 7268 24716 7296
rect 23658 7256 23664 7268
rect 23492 7228 23664 7256
rect 23201 7219 23259 7225
rect 23658 7216 23664 7228
rect 23716 7256 23722 7268
rect 24578 7256 24584 7268
rect 23716 7228 24584 7256
rect 23716 7216 23722 7228
rect 24578 7216 24584 7228
rect 24636 7216 24642 7268
rect 24670 7216 24676 7268
rect 24728 7256 24734 7268
rect 25516 7256 25544 7355
rect 24728 7228 25544 7256
rect 24728 7216 24734 7228
rect 21784 7160 22600 7188
rect 21784 7148 21790 7160
rect 1104 7098 32476 7120
rect 1104 7046 4871 7098
rect 4923 7046 4935 7098
rect 4987 7046 4999 7098
rect 5051 7046 5063 7098
rect 5115 7046 5127 7098
rect 5179 7046 12713 7098
rect 12765 7046 12777 7098
rect 12829 7046 12841 7098
rect 12893 7046 12905 7098
rect 12957 7046 12969 7098
rect 13021 7046 20555 7098
rect 20607 7046 20619 7098
rect 20671 7046 20683 7098
rect 20735 7046 20747 7098
rect 20799 7046 20811 7098
rect 20863 7046 28397 7098
rect 28449 7046 28461 7098
rect 28513 7046 28525 7098
rect 28577 7046 28589 7098
rect 28641 7046 28653 7098
rect 28705 7046 32476 7098
rect 1104 7024 32476 7046
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4246 6984 4252 6996
rect 4203 6956 4252 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 5261 6987 5319 6993
rect 5261 6953 5273 6987
rect 5307 6984 5319 6987
rect 5350 6984 5356 6996
rect 5307 6956 5356 6984
rect 5307 6953 5319 6956
rect 5261 6947 5319 6953
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5905 6987 5963 6993
rect 5905 6984 5917 6987
rect 5592 6956 5917 6984
rect 5592 6944 5598 6956
rect 5905 6953 5917 6956
rect 5951 6953 5963 6987
rect 5905 6947 5963 6953
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6420 6956 6561 6984
rect 6420 6944 6426 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 6549 6947 6607 6953
rect 13078 6944 13084 6996
rect 13136 6944 13142 6996
rect 16025 6987 16083 6993
rect 16025 6984 16037 6987
rect 15948 6956 16037 6984
rect 3050 6876 3056 6928
rect 3108 6876 3114 6928
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 3786 6848 3792 6860
rect 2639 6820 3792 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4264 6848 4292 6944
rect 12529 6919 12587 6925
rect 12176 6888 12388 6916
rect 4264 6820 4936 6848
rect 2682 6740 2688 6792
rect 2740 6789 2746 6792
rect 2740 6783 2789 6789
rect 2740 6749 2743 6783
rect 2777 6749 2789 6783
rect 2740 6743 2789 6749
rect 2740 6740 2746 6743
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3970 6780 3976 6792
rect 3384 6752 3976 6780
rect 3384 6740 3390 6752
rect 3970 6740 3976 6752
rect 4028 6780 4034 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 4028 6752 4077 6780
rect 4028 6740 4034 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4338 6780 4344 6792
rect 4295 6752 4344 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 4908 6789 4936 6820
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5040 6820 6040 6848
rect 5040 6808 5046 6820
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5316 6752 5733 6780
rect 5316 6740 5322 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 6012 6644 6040 6820
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 7708 6820 8432 6848
rect 7708 6808 7714 6820
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 7742 6780 7748 6792
rect 7607 6752 7748 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 8404 6789 8432 6820
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 8628 6820 9321 6848
rect 8628 6808 8634 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9398 6808 9404 6860
rect 9456 6808 9462 6860
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 9732 6820 10333 6848
rect 9732 6808 9738 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 12176 6848 12204 6888
rect 10321 6811 10379 6817
rect 11256 6820 12204 6848
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9548 6752 9781 6780
rect 9548 6740 9554 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 11256 6789 11284 6820
rect 12250 6808 12256 6860
rect 12308 6808 12314 6860
rect 12360 6848 12388 6888
rect 12529 6885 12541 6919
rect 12575 6885 12587 6919
rect 12529 6879 12587 6885
rect 12434 6848 12440 6860
rect 12360 6820 12440 6848
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 12544 6848 12572 6879
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 14369 6919 14427 6925
rect 14369 6916 14381 6919
rect 13872 6888 14381 6916
rect 13872 6876 13878 6888
rect 14369 6885 14381 6888
rect 14415 6885 14427 6919
rect 14369 6879 14427 6885
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 12544 6820 13277 6848
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 14737 6851 14795 6857
rect 14737 6817 14749 6851
rect 14783 6848 14795 6851
rect 14826 6848 14832 6860
rect 14783 6820 14832 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 14826 6808 14832 6820
rect 14884 6848 14890 6860
rect 15948 6848 15976 6956
rect 16025 6953 16037 6956
rect 16071 6953 16083 6987
rect 16025 6947 16083 6953
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 17405 6987 17463 6993
rect 17405 6984 17417 6987
rect 17276 6956 17417 6984
rect 17276 6944 17282 6956
rect 17405 6953 17417 6956
rect 17451 6953 17463 6987
rect 17405 6947 17463 6953
rect 17954 6944 17960 6996
rect 18012 6944 18018 6996
rect 20438 6944 20444 6996
rect 20496 6944 20502 6996
rect 22557 6987 22615 6993
rect 22557 6984 22569 6987
rect 22066 6956 22569 6984
rect 20806 6876 20812 6928
rect 20864 6916 20870 6928
rect 21358 6916 21364 6928
rect 20864 6888 21364 6916
rect 20864 6876 20870 6888
rect 21358 6876 21364 6888
rect 21416 6916 21422 6928
rect 21726 6916 21732 6928
rect 21416 6888 21732 6916
rect 21416 6876 21422 6888
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 16114 6848 16120 6860
rect 14884 6820 16120 6848
rect 14884 6808 14890 6820
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6848 17187 6851
rect 17310 6848 17316 6860
rect 17175 6820 17316 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 21913 6851 21971 6857
rect 17644 6820 19472 6848
rect 17644 6808 17650 6820
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 12158 6740 12164 6792
rect 12216 6740 12222 6792
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 12406 6752 13369 6780
rect 8573 6715 8631 6721
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 11057 6715 11115 6721
rect 8619 6684 9628 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 9600 6656 9628 6684
rect 11057 6681 11069 6715
rect 11103 6712 11115 6715
rect 12406 6712 12434 6752
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 15896 6752 15945 6780
rect 15896 6740 15902 6752
rect 15933 6749 15945 6752
rect 15979 6780 15991 6783
rect 16942 6780 16948 6792
rect 15979 6752 16948 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17034 6740 17040 6792
rect 17092 6740 17098 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 19444 6789 19472 6820
rect 20732 6820 21588 6848
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17276 6752 17877 6780
rect 17276 6740 17282 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19610 6780 19616 6792
rect 19475 6752 19616 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 18064 6712 18092 6743
rect 19610 6740 19616 6752
rect 19668 6780 19674 6792
rect 20346 6780 20352 6792
rect 19668 6752 20352 6780
rect 19668 6740 19674 6752
rect 20346 6740 20352 6752
rect 20404 6740 20410 6792
rect 20732 6789 20760 6820
rect 21560 6792 21588 6820
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 22066 6848 22094 6956
rect 22557 6953 22569 6956
rect 22603 6953 22615 6987
rect 22557 6947 22615 6953
rect 23845 6987 23903 6993
rect 23845 6953 23857 6987
rect 23891 6984 23903 6987
rect 24670 6984 24676 6996
rect 23891 6956 24676 6984
rect 23891 6953 23903 6956
rect 23845 6947 23903 6953
rect 24670 6944 24676 6956
rect 24728 6944 24734 6996
rect 22370 6876 22376 6928
rect 22428 6876 22434 6928
rect 21959 6820 22094 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 22554 6808 22560 6860
rect 22612 6848 22618 6860
rect 22612 6820 22968 6848
rect 22612 6808 22618 6820
rect 20625 6783 20683 6789
rect 20625 6749 20637 6783
rect 20671 6749 20683 6783
rect 20625 6743 20683 6749
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 11103 6684 12434 6712
rect 16408 6684 18092 6712
rect 20640 6712 20668 6743
rect 20898 6740 20904 6792
rect 20956 6740 20962 6792
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6780 21051 6783
rect 21082 6780 21088 6792
rect 21039 6752 21088 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 21450 6740 21456 6792
rect 21508 6740 21514 6792
rect 21542 6740 21548 6792
rect 21600 6740 21606 6792
rect 21726 6740 21732 6792
rect 21784 6740 21790 6792
rect 22525 6715 22583 6721
rect 22525 6712 22537 6715
rect 20640 6684 21864 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 6012 6616 9137 6644
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9582 6604 9588 6656
rect 9640 6604 9646 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 9766 6644 9772 6656
rect 9723 6616 9772 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 11425 6647 11483 6653
rect 11425 6613 11437 6647
rect 11471 6644 11483 6647
rect 11974 6644 11980 6656
rect 11471 6616 11980 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 16408 6653 16436 6684
rect 21836 6656 21864 6684
rect 22066 6684 22537 6712
rect 14277 6647 14335 6653
rect 14277 6644 14289 6647
rect 12492 6616 14289 6644
rect 12492 6604 12498 6616
rect 14277 6613 14289 6616
rect 14323 6613 14335 6647
rect 14277 6607 14335 6613
rect 16393 6647 16451 6653
rect 16393 6613 16405 6647
rect 16439 6613 16451 6647
rect 16393 6607 16451 6613
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 18196 6616 19625 6644
rect 18196 6604 18202 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 20070 6604 20076 6656
rect 20128 6644 20134 6656
rect 21082 6644 21088 6656
rect 20128 6616 21088 6644
rect 20128 6604 20134 6616
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 21818 6604 21824 6656
rect 21876 6644 21882 6656
rect 22066 6644 22094 6684
rect 22525 6681 22537 6684
rect 22571 6681 22583 6715
rect 22525 6675 22583 6681
rect 22741 6715 22799 6721
rect 22741 6681 22753 6715
rect 22787 6681 22799 6715
rect 22940 6712 22968 6820
rect 23014 6740 23020 6792
rect 23072 6780 23078 6792
rect 23661 6783 23719 6789
rect 23661 6780 23673 6783
rect 23072 6752 23673 6780
rect 23072 6740 23078 6752
rect 23661 6749 23673 6752
rect 23707 6749 23719 6783
rect 23661 6743 23719 6749
rect 23477 6715 23535 6721
rect 23477 6712 23489 6715
rect 22940 6684 23489 6712
rect 22741 6675 22799 6681
rect 23477 6681 23489 6684
rect 23523 6681 23535 6715
rect 23477 6675 23535 6681
rect 21876 6616 22094 6644
rect 22756 6644 22784 6675
rect 23290 6644 23296 6656
rect 22756 6616 23296 6644
rect 21876 6604 21882 6616
rect 23290 6604 23296 6616
rect 23348 6604 23354 6656
rect 1104 6554 32632 6576
rect 1104 6502 8792 6554
rect 8844 6502 8856 6554
rect 8908 6502 8920 6554
rect 8972 6502 8984 6554
rect 9036 6502 9048 6554
rect 9100 6502 16634 6554
rect 16686 6502 16698 6554
rect 16750 6502 16762 6554
rect 16814 6502 16826 6554
rect 16878 6502 16890 6554
rect 16942 6502 24476 6554
rect 24528 6502 24540 6554
rect 24592 6502 24604 6554
rect 24656 6502 24668 6554
rect 24720 6502 24732 6554
rect 24784 6502 32318 6554
rect 32370 6502 32382 6554
rect 32434 6502 32446 6554
rect 32498 6502 32510 6554
rect 32562 6502 32574 6554
rect 32626 6502 32632 6554
rect 1104 6480 32632 6502
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 4212 6412 4261 6440
rect 4212 6400 4218 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 9493 6443 9551 6449
rect 4672 6412 5120 6440
rect 4672 6400 4678 6412
rect 4338 6332 4344 6384
rect 4396 6372 4402 6384
rect 5092 6381 5120 6412
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 10134 6440 10140 6452
rect 9539 6412 10140 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 13722 6440 13728 6452
rect 13495 6412 13728 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6440 16911 6443
rect 17126 6440 17132 6452
rect 16899 6412 17132 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 21542 6400 21548 6452
rect 21600 6440 21606 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21600 6412 22017 6440
rect 21600 6400 21606 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 4893 6375 4951 6381
rect 4893 6372 4905 6375
rect 4396 6344 4905 6372
rect 4396 6332 4402 6344
rect 4893 6341 4905 6344
rect 4939 6341 4951 6375
rect 4893 6335 4951 6341
rect 5077 6375 5135 6381
rect 5077 6341 5089 6375
rect 5123 6341 5135 6375
rect 5077 6335 5135 6341
rect 5258 6332 5264 6384
rect 5316 6332 5322 6384
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6372 7987 6375
rect 7975 6344 9352 6372
rect 7975 6341 7987 6344
rect 7929 6335 7987 6341
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 4982 6304 4988 6316
rect 4488 6276 4988 6304
rect 4488 6264 4494 6276
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6304 8079 6307
rect 8294 6304 8300 6316
rect 8067 6276 8300 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 7852 6236 7880 6267
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8110 6236 8116 6248
rect 7852 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6236 8174 6248
rect 8496 6236 8524 6267
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9324 6313 9352 6344
rect 11514 6332 11520 6384
rect 11572 6372 11578 6384
rect 11572 6344 13216 6372
rect 11572 6332 11578 6344
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8628 6276 8677 6304
rect 8628 6264 8634 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 9490 6264 9496 6316
rect 9548 6264 9554 6316
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 12452 6276 13093 6304
rect 8168 6208 8524 6236
rect 8849 6239 8907 6245
rect 8168 6196 8174 6208
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 9508 6236 9536 6264
rect 12452 6245 12480 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13188 6248 13216 6344
rect 15672 6344 18460 6372
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 14826 6304 14832 6316
rect 14783 6276 14832 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 15672 6313 15700 6344
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16482 6304 16488 6316
rect 16172 6276 16488 6304
rect 16172 6264 16178 6276
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17310 6304 17316 6316
rect 17083 6276 17316 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17310 6264 17316 6276
rect 17368 6304 17374 6316
rect 18432 6313 18460 6344
rect 19610 6332 19616 6384
rect 19668 6332 19674 6384
rect 18417 6307 18475 6313
rect 17368 6276 18276 6304
rect 17368 6264 17374 6276
rect 8895 6208 9536 6236
rect 12437 6239 12495 6245
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 13170 6196 13176 6248
rect 13228 6196 13234 6248
rect 15856 6236 15884 6264
rect 15120 6208 15884 6236
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12434 6100 12440 6112
rect 12299 6072 12440 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 15120 6100 15148 6208
rect 17126 6196 17132 6248
rect 17184 6196 17190 6248
rect 17494 6196 17500 6248
rect 17552 6236 17558 6248
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17552 6208 17969 6236
rect 17552 6196 17558 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 15197 6171 15255 6177
rect 15197 6137 15209 6171
rect 15243 6168 15255 6171
rect 17218 6168 17224 6180
rect 15243 6140 17224 6168
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 17218 6128 17224 6140
rect 17276 6128 17282 6180
rect 15059 6072 15148 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16301 6103 16359 6109
rect 16301 6100 16313 6103
rect 16264 6072 16313 6100
rect 16264 6060 16270 6072
rect 16301 6069 16313 6072
rect 16347 6069 16359 6103
rect 16301 6063 16359 6069
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 18138 6100 18144 6112
rect 16540 6072 18144 6100
rect 16540 6060 16546 6072
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 18248 6100 18276 6276
rect 18417 6273 18429 6307
rect 18463 6304 18475 6307
rect 18598 6304 18604 6316
rect 18463 6276 18604 6304
rect 18463 6273 18475 6276
rect 18417 6267 18475 6273
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 19334 6128 19340 6180
rect 19392 6168 19398 6180
rect 19889 6171 19947 6177
rect 19889 6168 19901 6171
rect 19392 6140 19901 6168
rect 19392 6128 19398 6140
rect 19889 6137 19901 6140
rect 19935 6168 19947 6171
rect 20254 6168 20260 6180
rect 19935 6140 20260 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 20732 6168 20760 6267
rect 20806 6264 20812 6316
rect 20864 6264 20870 6316
rect 21082 6313 21088 6316
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 21058 6307 21088 6313
rect 21058 6273 21070 6307
rect 21058 6267 21088 6273
rect 20916 6236 20944 6267
rect 21082 6264 21088 6267
rect 21140 6264 21146 6316
rect 21174 6264 21180 6316
rect 21232 6264 21238 6316
rect 22462 6264 22468 6316
rect 22520 6264 22526 6316
rect 21450 6236 21456 6248
rect 20916 6208 21456 6236
rect 21450 6196 21456 6208
rect 21508 6236 21514 6248
rect 21726 6236 21732 6248
rect 21508 6208 21732 6236
rect 21508 6196 21514 6208
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 20898 6168 20904 6180
rect 20496 6140 20668 6168
rect 20732 6140 20904 6168
rect 20496 6128 20502 6140
rect 20533 6103 20591 6109
rect 20533 6100 20545 6103
rect 18248 6072 20545 6100
rect 20533 6069 20545 6072
rect 20579 6069 20591 6103
rect 20640 6100 20668 6140
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 22189 6103 22247 6109
rect 22189 6100 22201 6103
rect 20640 6072 22201 6100
rect 20533 6063 20591 6069
rect 22189 6069 22201 6072
rect 22235 6069 22247 6103
rect 22189 6063 22247 6069
rect 1104 6010 32476 6032
rect 1104 5958 4871 6010
rect 4923 5958 4935 6010
rect 4987 5958 4999 6010
rect 5051 5958 5063 6010
rect 5115 5958 5127 6010
rect 5179 5958 12713 6010
rect 12765 5958 12777 6010
rect 12829 5958 12841 6010
rect 12893 5958 12905 6010
rect 12957 5958 12969 6010
rect 13021 5958 20555 6010
rect 20607 5958 20619 6010
rect 20671 5958 20683 6010
rect 20735 5958 20747 6010
rect 20799 5958 20811 6010
rect 20863 5958 28397 6010
rect 28449 5958 28461 6010
rect 28513 5958 28525 6010
rect 28577 5958 28589 6010
rect 28641 5958 28653 6010
rect 28705 5958 32476 6010
rect 1104 5936 32476 5958
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12032 5868 12909 5896
rect 12032 5856 12038 5868
rect 12897 5865 12909 5868
rect 12943 5865 12955 5899
rect 12897 5859 12955 5865
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 13096 5828 13124 5859
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 16025 5899 16083 5905
rect 16025 5896 16037 5899
rect 13228 5868 16037 5896
rect 13228 5856 13234 5868
rect 16025 5865 16037 5868
rect 16071 5865 16083 5899
rect 16025 5859 16083 5865
rect 17126 5856 17132 5908
rect 17184 5856 17190 5908
rect 17497 5899 17555 5905
rect 17497 5865 17509 5899
rect 17543 5896 17555 5899
rect 18598 5896 18604 5908
rect 17543 5868 18604 5896
rect 17543 5865 17555 5868
rect 17497 5859 17555 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 20990 5896 20996 5908
rect 20763 5868 20996 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 21082 5856 21088 5908
rect 21140 5896 21146 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 21140 5868 21281 5896
rect 21140 5856 21146 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 21634 5856 21640 5908
rect 21692 5856 21698 5908
rect 22462 5856 22468 5908
rect 22520 5856 22526 5908
rect 13814 5828 13820 5840
rect 13096 5800 13820 5828
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 18138 5788 18144 5840
rect 18196 5828 18202 5840
rect 20438 5828 20444 5840
rect 18196 5800 20444 5828
rect 18196 5788 18202 5800
rect 20438 5788 20444 5800
rect 20496 5828 20502 5840
rect 20533 5831 20591 5837
rect 20533 5828 20545 5831
rect 20496 5800 20545 5828
rect 20496 5788 20502 5800
rect 20533 5797 20545 5800
rect 20579 5797 20591 5831
rect 20533 5791 20591 5797
rect 16206 5720 16212 5772
rect 16264 5720 16270 5772
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 17494 5760 17500 5772
rect 16347 5732 17500 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 20254 5720 20260 5772
rect 20312 5720 20318 5772
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12216 5664 13369 5692
rect 12216 5652 12222 5664
rect 13357 5661 13369 5664
rect 13403 5692 13415 5695
rect 14826 5692 14832 5704
rect 13403 5664 14832 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 17218 5692 17224 5704
rect 16715 5664 17224 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 17586 5652 17592 5704
rect 17644 5652 17650 5704
rect 21008 5692 21036 5856
rect 21542 5828 21548 5840
rect 21468 5800 21548 5828
rect 21082 5720 21088 5772
rect 21140 5760 21146 5772
rect 21468 5769 21496 5800
rect 21542 5788 21548 5800
rect 21600 5788 21606 5840
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 21140 5732 21465 5760
rect 21140 5720 21146 5732
rect 21453 5729 21465 5732
rect 21499 5729 21511 5763
rect 21453 5723 21511 5729
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 21008 5664 21189 5692
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21818 5692 21824 5704
rect 21591 5664 21824 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 22557 5695 22615 5701
rect 22557 5661 22569 5695
rect 22603 5692 22615 5695
rect 23014 5692 23020 5704
rect 22603 5664 23020 5692
rect 22603 5661 22615 5664
rect 22557 5655 22615 5661
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 17126 5624 17132 5636
rect 16500 5596 17132 5624
rect 16500 5565 16528 5596
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 16485 5559 16543 5565
rect 16485 5525 16497 5559
rect 16531 5525 16543 5559
rect 16485 5519 16543 5525
rect 16577 5559 16635 5565
rect 16577 5525 16589 5559
rect 16623 5556 16635 5559
rect 17310 5556 17316 5568
rect 16623 5528 17316 5556
rect 16623 5525 16635 5528
rect 16577 5519 16635 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 21726 5516 21732 5568
rect 21784 5556 21790 5568
rect 22097 5559 22155 5565
rect 22097 5556 22109 5559
rect 21784 5528 22109 5556
rect 21784 5516 21790 5528
rect 22097 5525 22109 5528
rect 22143 5525 22155 5559
rect 22097 5519 22155 5525
rect 1104 5466 32632 5488
rect 1104 5414 8792 5466
rect 8844 5414 8856 5466
rect 8908 5414 8920 5466
rect 8972 5414 8984 5466
rect 9036 5414 9048 5466
rect 9100 5414 16634 5466
rect 16686 5414 16698 5466
rect 16750 5414 16762 5466
rect 16814 5414 16826 5466
rect 16878 5414 16890 5466
rect 16942 5414 24476 5466
rect 24528 5414 24540 5466
rect 24592 5414 24604 5466
rect 24656 5414 24668 5466
rect 24720 5414 24732 5466
rect 24784 5414 32318 5466
rect 32370 5414 32382 5466
rect 32434 5414 32446 5466
rect 32498 5414 32510 5466
rect 32562 5414 32574 5466
rect 32626 5414 32632 5466
rect 1104 5392 32632 5414
rect 17034 5312 17040 5364
rect 17092 5312 17098 5364
rect 20625 5355 20683 5361
rect 20625 5321 20637 5355
rect 20671 5352 20683 5355
rect 20898 5352 20904 5364
rect 20671 5324 20904 5352
rect 20671 5321 20683 5324
rect 20625 5315 20683 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 21269 5355 21327 5361
rect 21269 5321 21281 5355
rect 21315 5352 21327 5355
rect 21818 5352 21824 5364
rect 21315 5324 21824 5352
rect 21315 5321 21327 5324
rect 21269 5315 21327 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 17126 5284 17132 5296
rect 16868 5256 17132 5284
rect 16868 5225 16896 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 21177 5287 21235 5293
rect 21177 5253 21189 5287
rect 21223 5284 21235 5287
rect 21726 5284 21732 5296
rect 21223 5256 21732 5284
rect 21223 5253 21235 5256
rect 21177 5247 21235 5253
rect 21726 5244 21732 5256
rect 21784 5244 21790 5296
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17494 5216 17500 5228
rect 17083 5188 17500 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17494 5176 17500 5188
rect 17552 5176 17558 5228
rect 19610 5176 19616 5228
rect 19668 5216 19674 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19668 5188 20177 5216
rect 19668 5176 19674 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 21082 5176 21088 5228
rect 21140 5176 21146 5228
rect 21358 5176 21364 5228
rect 21416 5176 21422 5228
rect 20254 4972 20260 5024
rect 20312 4972 20318 5024
rect 1104 4922 32476 4944
rect 1104 4870 4871 4922
rect 4923 4870 4935 4922
rect 4987 4870 4999 4922
rect 5051 4870 5063 4922
rect 5115 4870 5127 4922
rect 5179 4870 12713 4922
rect 12765 4870 12777 4922
rect 12829 4870 12841 4922
rect 12893 4870 12905 4922
rect 12957 4870 12969 4922
rect 13021 4870 20555 4922
rect 20607 4870 20619 4922
rect 20671 4870 20683 4922
rect 20735 4870 20747 4922
rect 20799 4870 20811 4922
rect 20863 4870 28397 4922
rect 28449 4870 28461 4922
rect 28513 4870 28525 4922
rect 28577 4870 28589 4922
rect 28641 4870 28653 4922
rect 28705 4870 32476 4922
rect 1104 4848 32476 4870
rect 1104 4378 32632 4400
rect 1104 4326 8792 4378
rect 8844 4326 8856 4378
rect 8908 4326 8920 4378
rect 8972 4326 8984 4378
rect 9036 4326 9048 4378
rect 9100 4326 16634 4378
rect 16686 4326 16698 4378
rect 16750 4326 16762 4378
rect 16814 4326 16826 4378
rect 16878 4326 16890 4378
rect 16942 4326 24476 4378
rect 24528 4326 24540 4378
rect 24592 4326 24604 4378
rect 24656 4326 24668 4378
rect 24720 4326 24732 4378
rect 24784 4326 32318 4378
rect 32370 4326 32382 4378
rect 32434 4326 32446 4378
rect 32498 4326 32510 4378
rect 32562 4326 32574 4378
rect 32626 4326 32632 4378
rect 1104 4304 32632 4326
rect 1104 3834 32476 3856
rect 1104 3782 4871 3834
rect 4923 3782 4935 3834
rect 4987 3782 4999 3834
rect 5051 3782 5063 3834
rect 5115 3782 5127 3834
rect 5179 3782 12713 3834
rect 12765 3782 12777 3834
rect 12829 3782 12841 3834
rect 12893 3782 12905 3834
rect 12957 3782 12969 3834
rect 13021 3782 20555 3834
rect 20607 3782 20619 3834
rect 20671 3782 20683 3834
rect 20735 3782 20747 3834
rect 20799 3782 20811 3834
rect 20863 3782 28397 3834
rect 28449 3782 28461 3834
rect 28513 3782 28525 3834
rect 28577 3782 28589 3834
rect 28641 3782 28653 3834
rect 28705 3782 32476 3834
rect 1104 3760 32476 3782
rect 1104 3290 32632 3312
rect 1104 3238 8792 3290
rect 8844 3238 8856 3290
rect 8908 3238 8920 3290
rect 8972 3238 8984 3290
rect 9036 3238 9048 3290
rect 9100 3238 16634 3290
rect 16686 3238 16698 3290
rect 16750 3238 16762 3290
rect 16814 3238 16826 3290
rect 16878 3238 16890 3290
rect 16942 3238 24476 3290
rect 24528 3238 24540 3290
rect 24592 3238 24604 3290
rect 24656 3238 24668 3290
rect 24720 3238 24732 3290
rect 24784 3238 32318 3290
rect 32370 3238 32382 3290
rect 32434 3238 32446 3290
rect 32498 3238 32510 3290
rect 32562 3238 32574 3290
rect 32626 3238 32632 3290
rect 1104 3216 32632 3238
rect 1104 2746 32476 2768
rect 1104 2694 4871 2746
rect 4923 2694 4935 2746
rect 4987 2694 4999 2746
rect 5051 2694 5063 2746
rect 5115 2694 5127 2746
rect 5179 2694 12713 2746
rect 12765 2694 12777 2746
rect 12829 2694 12841 2746
rect 12893 2694 12905 2746
rect 12957 2694 12969 2746
rect 13021 2694 20555 2746
rect 20607 2694 20619 2746
rect 20671 2694 20683 2746
rect 20735 2694 20747 2746
rect 20799 2694 20811 2746
rect 20863 2694 28397 2746
rect 28449 2694 28461 2746
rect 28513 2694 28525 2746
rect 28577 2694 28589 2746
rect 28641 2694 28653 2746
rect 28705 2694 32476 2746
rect 1104 2672 32476 2694
rect 1104 2202 32632 2224
rect 1104 2150 8792 2202
rect 8844 2150 8856 2202
rect 8908 2150 8920 2202
rect 8972 2150 8984 2202
rect 9036 2150 9048 2202
rect 9100 2150 16634 2202
rect 16686 2150 16698 2202
rect 16750 2150 16762 2202
rect 16814 2150 16826 2202
rect 16878 2150 16890 2202
rect 16942 2150 24476 2202
rect 24528 2150 24540 2202
rect 24592 2150 24604 2202
rect 24656 2150 24668 2202
rect 24720 2150 24732 2202
rect 24784 2150 32318 2202
rect 32370 2150 32382 2202
rect 32434 2150 32446 2202
rect 32498 2150 32510 2202
rect 32562 2150 32574 2202
rect 32626 2150 32632 2202
rect 1104 2128 32632 2150
rect 1104 1658 32476 1680
rect 1104 1606 4871 1658
rect 4923 1606 4935 1658
rect 4987 1606 4999 1658
rect 5051 1606 5063 1658
rect 5115 1606 5127 1658
rect 5179 1606 12713 1658
rect 12765 1606 12777 1658
rect 12829 1606 12841 1658
rect 12893 1606 12905 1658
rect 12957 1606 12969 1658
rect 13021 1606 20555 1658
rect 20607 1606 20619 1658
rect 20671 1606 20683 1658
rect 20735 1606 20747 1658
rect 20799 1606 20811 1658
rect 20863 1606 28397 1658
rect 28449 1606 28461 1658
rect 28513 1606 28525 1658
rect 28577 1606 28589 1658
rect 28641 1606 28653 1658
rect 28705 1606 32476 1658
rect 1104 1584 32476 1606
rect 1104 1114 32632 1136
rect 1104 1062 8792 1114
rect 8844 1062 8856 1114
rect 8908 1062 8920 1114
rect 8972 1062 8984 1114
rect 9036 1062 9048 1114
rect 9100 1062 16634 1114
rect 16686 1062 16698 1114
rect 16750 1062 16762 1114
rect 16814 1062 16826 1114
rect 16878 1062 16890 1114
rect 16942 1062 24476 1114
rect 24528 1062 24540 1114
rect 24592 1062 24604 1114
rect 24656 1062 24668 1114
rect 24720 1062 24732 1114
rect 24784 1062 32318 1114
rect 32370 1062 32382 1114
rect 32434 1062 32446 1114
rect 32498 1062 32510 1114
rect 32562 1062 32574 1114
rect 32626 1062 32632 1114
rect 1104 1040 32632 1062
<< via1 >>
rect 5356 20816 5408 20868
rect 10140 20816 10192 20868
rect 4896 20748 4948 20800
rect 15844 20748 15896 20800
rect 8792 20646 8844 20698
rect 8856 20646 8908 20698
rect 8920 20646 8972 20698
rect 8984 20646 9036 20698
rect 9048 20646 9100 20698
rect 16634 20646 16686 20698
rect 16698 20646 16750 20698
rect 16762 20646 16814 20698
rect 16826 20646 16878 20698
rect 16890 20646 16942 20698
rect 24476 20646 24528 20698
rect 24540 20646 24592 20698
rect 24604 20646 24656 20698
rect 24668 20646 24720 20698
rect 24732 20646 24784 20698
rect 32318 20646 32370 20698
rect 32382 20646 32434 20698
rect 32446 20646 32498 20698
rect 32510 20646 32562 20698
rect 32574 20646 32626 20698
rect 4436 20544 4488 20596
rect 4896 20587 4948 20596
rect 4896 20553 4905 20587
rect 4905 20553 4939 20587
rect 4939 20553 4948 20587
rect 4896 20544 4948 20553
rect 8116 20587 8168 20596
rect 8116 20553 8125 20587
rect 8125 20553 8159 20587
rect 8159 20553 8168 20587
rect 8116 20544 8168 20553
rect 9496 20587 9548 20596
rect 9496 20553 9505 20587
rect 9505 20553 9539 20587
rect 9539 20553 9548 20587
rect 9496 20544 9548 20553
rect 9680 20544 9732 20596
rect 13544 20587 13596 20596
rect 13544 20553 13553 20587
rect 13553 20553 13587 20587
rect 13587 20553 13596 20587
rect 13544 20544 13596 20553
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 17040 20587 17092 20596
rect 17040 20553 17049 20587
rect 17049 20553 17083 20587
rect 17083 20553 17092 20587
rect 17040 20544 17092 20553
rect 4804 20476 4856 20528
rect 11704 20519 11756 20528
rect 11704 20485 11713 20519
rect 11713 20485 11747 20519
rect 11747 20485 11756 20519
rect 11704 20476 11756 20485
rect 4712 20451 4764 20460
rect 4712 20417 4721 20451
rect 4721 20417 4755 20451
rect 4755 20417 4764 20451
rect 4712 20408 4764 20417
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 5540 20340 5592 20392
rect 6092 20272 6144 20324
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 10048 20408 10100 20460
rect 6828 20204 6880 20256
rect 9956 20272 10008 20324
rect 8116 20204 8168 20256
rect 10140 20383 10192 20392
rect 10140 20349 10149 20383
rect 10149 20349 10183 20383
rect 10183 20349 10192 20383
rect 10140 20340 10192 20349
rect 10784 20340 10836 20392
rect 10232 20272 10284 20324
rect 10968 20408 11020 20460
rect 15384 20476 15436 20528
rect 11980 20451 12032 20460
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 13636 20408 13688 20460
rect 13820 20272 13872 20324
rect 15384 20340 15436 20392
rect 17408 20476 17460 20528
rect 16396 20408 16448 20460
rect 18604 20408 18656 20460
rect 18972 20408 19024 20460
rect 20168 20408 20220 20460
rect 20260 20408 20312 20460
rect 20904 20408 20956 20460
rect 23572 20408 23624 20460
rect 26240 20408 26292 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27804 20451 27856 20460
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 30472 20408 30524 20460
rect 17500 20340 17552 20392
rect 17408 20272 17460 20324
rect 22100 20340 22152 20392
rect 25964 20340 26016 20392
rect 15752 20204 15804 20256
rect 23020 20272 23072 20324
rect 18880 20204 18932 20256
rect 20444 20204 20496 20256
rect 24952 20204 25004 20256
rect 29184 20247 29236 20256
rect 29184 20213 29193 20247
rect 29193 20213 29227 20247
rect 29227 20213 29236 20247
rect 29184 20204 29236 20213
rect 29736 20383 29788 20392
rect 29736 20349 29745 20383
rect 29745 20349 29779 20383
rect 29779 20349 29788 20383
rect 29736 20340 29788 20349
rect 31668 20247 31720 20256
rect 31668 20213 31677 20247
rect 31677 20213 31711 20247
rect 31711 20213 31720 20247
rect 31668 20204 31720 20213
rect 4871 20102 4923 20154
rect 4935 20102 4987 20154
rect 4999 20102 5051 20154
rect 5063 20102 5115 20154
rect 5127 20102 5179 20154
rect 12713 20102 12765 20154
rect 12777 20102 12829 20154
rect 12841 20102 12893 20154
rect 12905 20102 12957 20154
rect 12969 20102 13021 20154
rect 20555 20102 20607 20154
rect 20619 20102 20671 20154
rect 20683 20102 20735 20154
rect 20747 20102 20799 20154
rect 20811 20102 20863 20154
rect 28397 20102 28449 20154
rect 28461 20102 28513 20154
rect 28525 20102 28577 20154
rect 28589 20102 28641 20154
rect 28653 20102 28705 20154
rect 4712 20000 4764 20052
rect 5356 20043 5408 20052
rect 5356 20009 5365 20043
rect 5365 20009 5399 20043
rect 5399 20009 5408 20043
rect 5356 20000 5408 20009
rect 6000 20000 6052 20052
rect 8208 20000 8260 20052
rect 8576 19932 8628 19984
rect 14188 20000 14240 20052
rect 15016 20000 15068 20052
rect 2964 19864 3016 19916
rect 8208 19864 8260 19916
rect 3240 19839 3292 19848
rect 3240 19805 3249 19839
rect 3249 19805 3283 19839
rect 3283 19805 3292 19839
rect 3240 19796 3292 19805
rect 4068 19796 4120 19848
rect 7012 19796 7064 19848
rect 8116 19796 8168 19848
rect 15292 19864 15344 19916
rect 18972 20000 19024 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20444 20000 20496 20052
rect 22100 20043 22152 20052
rect 22100 20009 22109 20043
rect 22109 20009 22143 20043
rect 22143 20009 22152 20043
rect 22100 20000 22152 20009
rect 27804 20000 27856 20052
rect 20996 19932 21048 19984
rect 2780 19703 2832 19712
rect 2780 19669 2789 19703
rect 2789 19669 2823 19703
rect 2823 19669 2832 19703
rect 2780 19660 2832 19669
rect 3516 19728 3568 19780
rect 4344 19660 4396 19712
rect 8208 19728 8260 19780
rect 11244 19796 11296 19848
rect 9680 19728 9732 19780
rect 12164 19796 12216 19848
rect 12624 19796 12676 19848
rect 13728 19839 13780 19848
rect 13728 19805 13737 19839
rect 13737 19805 13771 19839
rect 13771 19805 13780 19839
rect 13728 19796 13780 19805
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 15384 19796 15436 19848
rect 12072 19728 12124 19780
rect 8484 19703 8536 19712
rect 8484 19669 8493 19703
rect 8493 19669 8527 19703
rect 8527 19669 8536 19703
rect 8484 19660 8536 19669
rect 9312 19660 9364 19712
rect 9588 19660 9640 19712
rect 10968 19660 11020 19712
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 13544 19660 13596 19712
rect 14648 19728 14700 19780
rect 17408 19796 17460 19848
rect 18696 19796 18748 19848
rect 19800 19796 19852 19848
rect 19984 19839 20036 19848
rect 19984 19805 20017 19839
rect 20017 19805 20036 19839
rect 22376 19864 22428 19916
rect 24860 19907 24912 19916
rect 24860 19873 24869 19907
rect 24869 19873 24903 19907
rect 24903 19873 24912 19907
rect 24860 19864 24912 19873
rect 19984 19796 20036 19805
rect 15752 19771 15804 19780
rect 15752 19737 15786 19771
rect 15786 19737 15804 19771
rect 15752 19728 15804 19737
rect 18604 19728 18656 19780
rect 20076 19728 20128 19780
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 22284 19796 22336 19848
rect 23020 19839 23072 19848
rect 23020 19805 23029 19839
rect 23029 19805 23063 19839
rect 23063 19805 23072 19839
rect 23020 19796 23072 19805
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 29460 19932 29512 19984
rect 26792 19907 26844 19916
rect 26792 19873 26801 19907
rect 26801 19873 26835 19907
rect 26835 19873 26844 19907
rect 26792 19864 26844 19873
rect 26700 19839 26752 19848
rect 26700 19805 26709 19839
rect 26709 19805 26743 19839
rect 26743 19805 26752 19839
rect 26700 19796 26752 19805
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 28356 19796 28408 19848
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 30288 19796 30340 19848
rect 30932 19796 30984 19848
rect 31944 19796 31996 19848
rect 17040 19660 17092 19712
rect 18788 19660 18840 19712
rect 19984 19660 20036 19712
rect 20904 19660 20956 19712
rect 25964 19660 26016 19712
rect 27896 19703 27948 19712
rect 27896 19669 27905 19703
rect 27905 19669 27939 19703
rect 27939 19669 27948 19703
rect 27896 19660 27948 19669
rect 31576 19660 31628 19712
rect 8792 19558 8844 19610
rect 8856 19558 8908 19610
rect 8920 19558 8972 19610
rect 8984 19558 9036 19610
rect 9048 19558 9100 19610
rect 16634 19558 16686 19610
rect 16698 19558 16750 19610
rect 16762 19558 16814 19610
rect 16826 19558 16878 19610
rect 16890 19558 16942 19610
rect 24476 19558 24528 19610
rect 24540 19558 24592 19610
rect 24604 19558 24656 19610
rect 24668 19558 24720 19610
rect 24732 19558 24784 19610
rect 32318 19558 32370 19610
rect 32382 19558 32434 19610
rect 32446 19558 32498 19610
rect 32510 19558 32562 19610
rect 32574 19558 32626 19610
rect 1768 19499 1820 19508
rect 1768 19465 1777 19499
rect 1777 19465 1811 19499
rect 1811 19465 1820 19499
rect 1768 19456 1820 19465
rect 3516 19456 3568 19508
rect 6552 19456 6604 19508
rect 9680 19456 9732 19508
rect 12164 19456 12216 19508
rect 2780 19388 2832 19440
rect 9036 19388 9088 19440
rect 9220 19388 9272 19440
rect 9496 19431 9548 19440
rect 9496 19397 9505 19431
rect 9505 19397 9539 19431
rect 9539 19397 9548 19431
rect 9496 19388 9548 19397
rect 10048 19388 10100 19440
rect 11152 19388 11204 19440
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 3148 19320 3200 19372
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 2964 19252 3016 19304
rect 3424 19320 3476 19372
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 7104 19320 7156 19372
rect 3976 19252 4028 19304
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 8024 19320 8076 19372
rect 8208 19320 8260 19372
rect 8576 19320 8628 19372
rect 9588 19320 9640 19372
rect 9956 19320 10008 19372
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 16396 19456 16448 19508
rect 17132 19456 17184 19508
rect 18604 19499 18656 19508
rect 18604 19465 18613 19499
rect 18613 19465 18647 19499
rect 18647 19465 18656 19499
rect 18604 19456 18656 19465
rect 20904 19456 20956 19508
rect 20996 19456 21048 19508
rect 26700 19456 26752 19508
rect 26792 19456 26844 19508
rect 28356 19499 28408 19508
rect 28356 19465 28365 19499
rect 28365 19465 28399 19499
rect 28399 19465 28408 19499
rect 28356 19456 28408 19465
rect 29184 19456 29236 19508
rect 13084 19388 13136 19440
rect 15292 19388 15344 19440
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 13452 19320 13504 19372
rect 14648 19363 14700 19372
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 16488 19320 16540 19372
rect 17040 19320 17092 19372
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 19524 19320 19576 19372
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 20444 19320 20496 19372
rect 22192 19388 22244 19440
rect 5816 19184 5868 19236
rect 8024 19184 8076 19236
rect 9588 19184 9640 19236
rect 14464 19184 14516 19236
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 7196 19116 7248 19168
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 9036 19116 9088 19168
rect 9404 19116 9456 19168
rect 14556 19116 14608 19168
rect 20168 19252 20220 19304
rect 22100 19320 22152 19372
rect 21180 19252 21232 19304
rect 22008 19252 22060 19304
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 23204 19363 23256 19372
rect 23204 19329 23213 19363
rect 23213 19329 23247 19363
rect 23247 19329 23256 19363
rect 23204 19320 23256 19329
rect 25872 19388 25924 19440
rect 22744 19252 22796 19304
rect 18696 19184 18748 19236
rect 26240 19320 26292 19372
rect 27436 19388 27488 19440
rect 28816 19388 28868 19440
rect 31484 19456 31536 19508
rect 26516 19320 26568 19372
rect 27896 19320 27948 19372
rect 25964 19252 26016 19304
rect 26424 19252 26476 19304
rect 24860 19184 24912 19236
rect 25872 19227 25924 19236
rect 25872 19193 25881 19227
rect 25881 19193 25915 19227
rect 25915 19193 25924 19227
rect 25872 19184 25924 19193
rect 15844 19116 15896 19168
rect 17132 19116 17184 19168
rect 18420 19116 18472 19168
rect 19708 19116 19760 19168
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 22652 19116 22704 19168
rect 26332 19116 26384 19168
rect 27344 19116 27396 19168
rect 4871 19014 4923 19066
rect 4935 19014 4987 19066
rect 4999 19014 5051 19066
rect 5063 19014 5115 19066
rect 5127 19014 5179 19066
rect 12713 19014 12765 19066
rect 12777 19014 12829 19066
rect 12841 19014 12893 19066
rect 12905 19014 12957 19066
rect 12969 19014 13021 19066
rect 20555 19014 20607 19066
rect 20619 19014 20671 19066
rect 20683 19014 20735 19066
rect 20747 19014 20799 19066
rect 20811 19014 20863 19066
rect 28397 19014 28449 19066
rect 28461 19014 28513 19066
rect 28525 19014 28577 19066
rect 28589 19014 28641 19066
rect 28653 19014 28705 19066
rect 2596 18912 2648 18964
rect 4344 18912 4396 18964
rect 7104 18912 7156 18964
rect 2228 18844 2280 18896
rect 4068 18844 4120 18896
rect 5816 18776 5868 18828
rect 8484 18912 8536 18964
rect 8668 18912 8720 18964
rect 9496 18912 9548 18964
rect 10876 18912 10928 18964
rect 11060 18844 11112 18896
rect 11888 18844 11940 18896
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 2964 18708 3016 18760
rect 3424 18708 3476 18760
rect 10600 18776 10652 18828
rect 14556 18912 14608 18964
rect 17408 18912 17460 18964
rect 18696 18955 18748 18964
rect 18696 18921 18705 18955
rect 18705 18921 18739 18955
rect 18739 18921 18748 18955
rect 18696 18912 18748 18921
rect 20260 18912 20312 18964
rect 21180 18955 21232 18964
rect 21180 18921 21189 18955
rect 21189 18921 21223 18955
rect 21223 18921 21232 18955
rect 21180 18912 21232 18921
rect 21272 18912 21324 18964
rect 13452 18844 13504 18896
rect 2228 18615 2280 18624
rect 2228 18581 2237 18615
rect 2237 18581 2271 18615
rect 2271 18581 2280 18615
rect 2228 18572 2280 18581
rect 2872 18572 2924 18624
rect 4068 18572 4120 18624
rect 8116 18708 8168 18760
rect 8300 18708 8352 18760
rect 7104 18572 7156 18624
rect 8668 18640 8720 18692
rect 9312 18708 9364 18760
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9680 18708 9732 18760
rect 10416 18708 10468 18760
rect 11060 18708 11112 18760
rect 14740 18776 14792 18828
rect 19616 18844 19668 18896
rect 19708 18887 19760 18896
rect 19708 18853 19717 18887
rect 19717 18853 19751 18887
rect 19751 18853 19760 18887
rect 19708 18844 19760 18853
rect 19800 18844 19852 18896
rect 9404 18572 9456 18624
rect 9956 18572 10008 18624
rect 11152 18683 11204 18692
rect 11152 18649 11161 18683
rect 11161 18649 11195 18683
rect 11195 18649 11204 18683
rect 11152 18640 11204 18649
rect 11336 18572 11388 18624
rect 12532 18708 12584 18760
rect 13268 18708 13320 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13084 18640 13136 18692
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 15476 18708 15528 18760
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 15936 18708 15988 18760
rect 15568 18640 15620 18692
rect 12440 18572 12492 18624
rect 12716 18572 12768 18624
rect 14464 18572 14516 18624
rect 15844 18572 15896 18624
rect 16304 18572 16356 18624
rect 16488 18615 16540 18624
rect 16488 18581 16497 18615
rect 16497 18581 16531 18615
rect 16531 18581 16540 18615
rect 16488 18572 16540 18581
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 18880 18819 18932 18828
rect 18880 18785 18889 18819
rect 18889 18785 18923 18819
rect 18923 18785 18932 18819
rect 18880 18776 18932 18785
rect 22376 18887 22428 18896
rect 22376 18853 22385 18887
rect 22385 18853 22419 18887
rect 22419 18853 22428 18887
rect 22376 18844 22428 18853
rect 23572 18887 23624 18896
rect 23572 18853 23581 18887
rect 23581 18853 23615 18887
rect 23615 18853 23624 18887
rect 23572 18844 23624 18853
rect 26516 18955 26568 18964
rect 26516 18921 26525 18955
rect 26525 18921 26559 18955
rect 26559 18921 26568 18955
rect 26516 18912 26568 18921
rect 27436 18912 27488 18964
rect 28080 18955 28132 18964
rect 28080 18921 28089 18955
rect 28089 18921 28123 18955
rect 28123 18921 28132 18955
rect 28080 18912 28132 18921
rect 30472 18912 30524 18964
rect 26240 18844 26292 18896
rect 18512 18708 18564 18760
rect 20444 18708 20496 18760
rect 19524 18640 19576 18692
rect 20352 18640 20404 18692
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 18880 18572 18932 18624
rect 21272 18708 21324 18760
rect 22008 18751 22060 18760
rect 22008 18717 22017 18751
rect 22017 18717 22051 18751
rect 22051 18717 22060 18751
rect 22008 18708 22060 18717
rect 23204 18708 23256 18760
rect 21456 18640 21508 18692
rect 24400 18708 24452 18760
rect 25136 18708 25188 18760
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 27344 18708 27396 18760
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 28724 18708 28776 18760
rect 24860 18640 24912 18692
rect 31576 18708 31628 18760
rect 30288 18640 30340 18692
rect 30932 18683 30984 18692
rect 30932 18649 30950 18683
rect 30950 18649 30984 18683
rect 30932 18640 30984 18649
rect 23388 18615 23440 18624
rect 23388 18581 23397 18615
rect 23397 18581 23431 18615
rect 23431 18581 23440 18615
rect 23388 18572 23440 18581
rect 25964 18572 26016 18624
rect 29184 18572 29236 18624
rect 32036 18572 32088 18624
rect 8792 18470 8844 18522
rect 8856 18470 8908 18522
rect 8920 18470 8972 18522
rect 8984 18470 9036 18522
rect 9048 18470 9100 18522
rect 16634 18470 16686 18522
rect 16698 18470 16750 18522
rect 16762 18470 16814 18522
rect 16826 18470 16878 18522
rect 16890 18470 16942 18522
rect 24476 18470 24528 18522
rect 24540 18470 24592 18522
rect 24604 18470 24656 18522
rect 24668 18470 24720 18522
rect 24732 18470 24784 18522
rect 32318 18470 32370 18522
rect 32382 18470 32434 18522
rect 32446 18470 32498 18522
rect 32510 18470 32562 18522
rect 32574 18470 32626 18522
rect 2596 18411 2648 18420
rect 2596 18377 2605 18411
rect 2605 18377 2639 18411
rect 2639 18377 2648 18411
rect 2596 18368 2648 18377
rect 3240 18368 3292 18420
rect 6920 18368 6972 18420
rect 8484 18368 8536 18420
rect 9404 18368 9456 18420
rect 10416 18368 10468 18420
rect 12624 18368 12676 18420
rect 2412 18300 2464 18352
rect 2688 18164 2740 18216
rect 3056 18275 3108 18284
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 5356 18300 5408 18352
rect 7288 18300 7340 18352
rect 8392 18300 8444 18352
rect 4436 18275 4488 18284
rect 4436 18241 4470 18275
rect 4470 18241 4488 18275
rect 4436 18232 4488 18241
rect 8024 18232 8076 18284
rect 9956 18343 10008 18352
rect 9956 18309 9965 18343
rect 9965 18309 9999 18343
rect 9999 18309 10008 18343
rect 9956 18300 10008 18309
rect 13636 18368 13688 18420
rect 15476 18368 15528 18420
rect 18420 18368 18472 18420
rect 18512 18368 18564 18420
rect 19616 18368 19668 18420
rect 20260 18368 20312 18420
rect 20352 18368 20404 18420
rect 20996 18368 21048 18420
rect 21456 18368 21508 18420
rect 22100 18411 22152 18420
rect 22100 18377 22109 18411
rect 22109 18377 22143 18411
rect 22143 18377 22152 18411
rect 22100 18368 22152 18377
rect 22744 18411 22796 18420
rect 22744 18377 22753 18411
rect 22753 18377 22787 18411
rect 22787 18377 22796 18411
rect 22744 18368 22796 18377
rect 23388 18368 23440 18420
rect 26424 18411 26476 18420
rect 26424 18377 26433 18411
rect 26433 18377 26467 18411
rect 26467 18377 26476 18411
rect 26424 18368 26476 18377
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 7104 18164 7156 18216
rect 7656 18164 7708 18216
rect 9680 18232 9732 18284
rect 11060 18275 11112 18284
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 11428 18232 11480 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 12900 18232 12952 18284
rect 18788 18300 18840 18352
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 14924 18232 14976 18284
rect 15660 18232 15712 18284
rect 7012 18139 7064 18148
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 8576 18096 8628 18148
rect 8668 18096 8720 18148
rect 2136 18028 2188 18080
rect 2228 18028 2280 18080
rect 6092 18028 6144 18080
rect 7196 18071 7248 18080
rect 7196 18037 7205 18071
rect 7205 18037 7239 18071
rect 7239 18037 7248 18071
rect 7196 18028 7248 18037
rect 7564 18028 7616 18080
rect 8024 18028 8076 18080
rect 12900 18096 12952 18148
rect 15476 18164 15528 18216
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 15936 18232 15988 18284
rect 20904 18300 20956 18352
rect 20260 18232 20312 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 22100 18232 22152 18284
rect 22560 18232 22612 18284
rect 31668 18300 31720 18352
rect 22744 18232 22796 18284
rect 24032 18275 24084 18284
rect 24032 18241 24041 18275
rect 24041 18241 24075 18275
rect 24075 18241 24084 18275
rect 24032 18232 24084 18241
rect 24400 18232 24452 18284
rect 24860 18232 24912 18284
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 26332 18232 26384 18284
rect 27436 18275 27488 18284
rect 27436 18241 27445 18275
rect 27445 18241 27479 18275
rect 27479 18241 27488 18275
rect 27436 18232 27488 18241
rect 29184 18232 29236 18284
rect 19248 18207 19300 18216
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 15016 18139 15068 18148
rect 15016 18105 15025 18139
rect 15025 18105 15059 18139
rect 15059 18105 15068 18139
rect 15016 18096 15068 18105
rect 18788 18096 18840 18148
rect 29092 18207 29144 18216
rect 29092 18173 29101 18207
rect 29101 18173 29135 18207
rect 29135 18173 29144 18207
rect 29092 18164 29144 18173
rect 19524 18139 19576 18148
rect 19524 18105 19533 18139
rect 19533 18105 19567 18139
rect 19567 18105 19576 18139
rect 19524 18096 19576 18105
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 11704 18028 11756 18080
rect 12440 18028 12492 18080
rect 13728 18028 13780 18080
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 14372 18028 14424 18080
rect 15292 18028 15344 18080
rect 15384 18028 15436 18080
rect 15660 18028 15712 18080
rect 15936 18028 15988 18080
rect 16120 18028 16172 18080
rect 17408 18028 17460 18080
rect 22008 18096 22060 18148
rect 19708 18071 19760 18080
rect 19708 18037 19717 18071
rect 19717 18037 19751 18071
rect 19751 18037 19760 18071
rect 19708 18028 19760 18037
rect 20168 18028 20220 18080
rect 23388 18028 23440 18080
rect 25228 18028 25280 18080
rect 27252 18071 27304 18080
rect 27252 18037 27261 18071
rect 27261 18037 27295 18071
rect 27295 18037 27304 18071
rect 27252 18028 27304 18037
rect 30380 18028 30432 18080
rect 31576 18071 31628 18080
rect 31576 18037 31585 18071
rect 31585 18037 31619 18071
rect 31619 18037 31628 18071
rect 31576 18028 31628 18037
rect 4871 17926 4923 17978
rect 4935 17926 4987 17978
rect 4999 17926 5051 17978
rect 5063 17926 5115 17978
rect 5127 17926 5179 17978
rect 12713 17926 12765 17978
rect 12777 17926 12829 17978
rect 12841 17926 12893 17978
rect 12905 17926 12957 17978
rect 12969 17926 13021 17978
rect 20555 17926 20607 17978
rect 20619 17926 20671 17978
rect 20683 17926 20735 17978
rect 20747 17926 20799 17978
rect 20811 17926 20863 17978
rect 28397 17926 28449 17978
rect 28461 17926 28513 17978
rect 28525 17926 28577 17978
rect 28589 17926 28641 17978
rect 28653 17926 28705 17978
rect 2412 17824 2464 17876
rect 3056 17824 3108 17876
rect 3608 17824 3660 17876
rect 3976 17824 4028 17876
rect 3424 17756 3476 17808
rect 4436 17867 4488 17876
rect 4436 17833 4445 17867
rect 4445 17833 4479 17867
rect 4479 17833 4488 17867
rect 4436 17824 4488 17833
rect 3148 17688 3200 17740
rect 3056 17620 3108 17672
rect 2136 17595 2188 17604
rect 2136 17561 2145 17595
rect 2145 17561 2179 17595
rect 2179 17561 2188 17595
rect 2136 17552 2188 17561
rect 2044 17484 2096 17536
rect 3148 17552 3200 17604
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 6092 17595 6144 17604
rect 6092 17561 6101 17595
rect 6101 17561 6135 17595
rect 6135 17561 6144 17595
rect 6092 17552 6144 17561
rect 3792 17484 3844 17536
rect 5356 17527 5408 17536
rect 5356 17493 5365 17527
rect 5365 17493 5399 17527
rect 5399 17493 5408 17527
rect 5356 17484 5408 17493
rect 10048 17824 10100 17876
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 11980 17824 12032 17876
rect 8024 17756 8076 17808
rect 8300 17756 8352 17808
rect 10232 17756 10284 17808
rect 10600 17799 10652 17808
rect 10600 17765 10609 17799
rect 10609 17765 10643 17799
rect 10643 17765 10652 17799
rect 10600 17756 10652 17765
rect 8392 17620 8444 17672
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 9864 17620 9916 17672
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 11152 17756 11204 17808
rect 11704 17799 11756 17808
rect 11704 17765 11713 17799
rect 11713 17765 11747 17799
rect 11747 17765 11756 17799
rect 11704 17756 11756 17765
rect 14740 17824 14792 17876
rect 11152 17620 11204 17672
rect 6736 17552 6788 17604
rect 7564 17595 7616 17604
rect 7564 17561 7573 17595
rect 7573 17561 7607 17595
rect 7607 17561 7616 17595
rect 7564 17552 7616 17561
rect 7748 17595 7800 17604
rect 7748 17561 7757 17595
rect 7757 17561 7791 17595
rect 7791 17561 7800 17595
rect 7748 17552 7800 17561
rect 11060 17552 11112 17604
rect 11336 17620 11388 17672
rect 12716 17756 12768 17808
rect 14372 17756 14424 17808
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 12440 17595 12492 17604
rect 12440 17561 12449 17595
rect 12449 17561 12483 17595
rect 12483 17561 12492 17595
rect 12440 17552 12492 17561
rect 12532 17595 12584 17604
rect 12532 17561 12541 17595
rect 12541 17561 12575 17595
rect 12575 17561 12584 17595
rect 12532 17552 12584 17561
rect 13452 17620 13504 17672
rect 14280 17620 14332 17672
rect 15200 17824 15252 17876
rect 15292 17824 15344 17876
rect 19524 17824 19576 17876
rect 19892 17824 19944 17876
rect 23204 17824 23256 17876
rect 23756 17824 23808 17876
rect 25136 17824 25188 17876
rect 31116 17824 31168 17876
rect 19432 17756 19484 17808
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 15384 17620 15436 17672
rect 16212 17731 16264 17740
rect 16212 17697 16221 17731
rect 16221 17697 16255 17731
rect 16255 17697 16264 17731
rect 16212 17688 16264 17697
rect 8300 17484 8352 17536
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 11980 17484 12032 17536
rect 12900 17552 12952 17604
rect 13176 17552 13228 17604
rect 13268 17552 13320 17604
rect 13728 17595 13780 17604
rect 13728 17561 13737 17595
rect 13737 17561 13771 17595
rect 13771 17561 13780 17595
rect 13728 17552 13780 17561
rect 12716 17484 12768 17536
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 17776 17688 17828 17740
rect 19708 17756 19760 17808
rect 20904 17756 20956 17808
rect 23572 17756 23624 17808
rect 17132 17552 17184 17604
rect 17408 17620 17460 17672
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 17684 17484 17736 17536
rect 18420 17663 18472 17672
rect 18420 17629 18426 17663
rect 18426 17629 18460 17663
rect 18460 17629 18472 17663
rect 18420 17620 18472 17629
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 18880 17663 18932 17672
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 21088 17688 21140 17740
rect 23112 17688 23164 17740
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 20260 17620 20312 17672
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 24860 17620 24912 17672
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 19248 17552 19300 17604
rect 20720 17552 20772 17604
rect 21088 17552 21140 17604
rect 23480 17552 23532 17604
rect 23664 17552 23716 17604
rect 19340 17484 19392 17536
rect 19984 17484 20036 17536
rect 23296 17484 23348 17536
rect 24308 17484 24360 17536
rect 24952 17595 25004 17604
rect 24952 17561 24961 17595
rect 24961 17561 24995 17595
rect 24995 17561 25004 17595
rect 24952 17552 25004 17561
rect 26608 17552 26660 17604
rect 28724 17620 28776 17672
rect 30288 17620 30340 17672
rect 31852 17620 31904 17672
rect 29736 17552 29788 17604
rect 31576 17552 31628 17604
rect 25780 17484 25832 17536
rect 26240 17484 26292 17536
rect 27436 17484 27488 17536
rect 29828 17484 29880 17536
rect 29920 17527 29972 17536
rect 29920 17493 29929 17527
rect 29929 17493 29963 17527
rect 29963 17493 29972 17527
rect 29920 17484 29972 17493
rect 30012 17484 30064 17536
rect 31852 17484 31904 17536
rect 8792 17382 8844 17434
rect 8856 17382 8908 17434
rect 8920 17382 8972 17434
rect 8984 17382 9036 17434
rect 9048 17382 9100 17434
rect 16634 17382 16686 17434
rect 16698 17382 16750 17434
rect 16762 17382 16814 17434
rect 16826 17382 16878 17434
rect 16890 17382 16942 17434
rect 24476 17382 24528 17434
rect 24540 17382 24592 17434
rect 24604 17382 24656 17434
rect 24668 17382 24720 17434
rect 24732 17382 24784 17434
rect 32318 17382 32370 17434
rect 32382 17382 32434 17434
rect 32446 17382 32498 17434
rect 32510 17382 32562 17434
rect 32574 17382 32626 17434
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 3424 17280 3476 17332
rect 3608 17280 3660 17332
rect 3056 17212 3108 17264
rect 2688 17144 2740 17196
rect 3240 17144 3292 17196
rect 4160 17144 4212 17196
rect 4344 17187 4396 17196
rect 4344 17153 4378 17187
rect 4378 17153 4396 17187
rect 4344 17144 4396 17153
rect 5540 17280 5592 17332
rect 8208 17280 8260 17332
rect 7012 17212 7064 17264
rect 9128 17212 9180 17264
rect 9864 17280 9916 17332
rect 9680 17212 9732 17264
rect 9956 17212 10008 17264
rect 10140 17212 10192 17264
rect 6000 17144 6052 17196
rect 6092 17144 6144 17196
rect 9864 17144 9916 17196
rect 11244 17212 11296 17264
rect 11796 17212 11848 17264
rect 12532 17280 12584 17332
rect 12716 17323 12768 17332
rect 12716 17289 12725 17323
rect 12725 17289 12759 17323
rect 12759 17289 12768 17323
rect 12716 17280 12768 17289
rect 12900 17323 12952 17332
rect 12900 17289 12909 17323
rect 12909 17289 12943 17323
rect 12943 17289 12952 17323
rect 12900 17280 12952 17289
rect 16488 17280 16540 17332
rect 17132 17280 17184 17332
rect 19524 17280 19576 17332
rect 19800 17323 19852 17332
rect 19800 17289 19809 17323
rect 19809 17289 19843 17323
rect 19843 17289 19852 17323
rect 19800 17280 19852 17289
rect 20260 17323 20312 17332
rect 20260 17289 20269 17323
rect 20269 17289 20303 17323
rect 20303 17289 20312 17323
rect 20260 17280 20312 17289
rect 23480 17280 23532 17332
rect 26056 17280 26108 17332
rect 3332 17008 3384 17060
rect 2044 16940 2096 16992
rect 3056 16940 3108 16992
rect 3424 16940 3476 16992
rect 7104 17119 7156 17128
rect 7104 17085 7113 17119
rect 7113 17085 7147 17119
rect 7147 17085 7156 17119
rect 7104 17076 7156 17085
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 8116 17119 8168 17128
rect 8116 17085 8125 17119
rect 8125 17085 8159 17119
rect 8159 17085 8168 17119
rect 8116 17076 8168 17085
rect 9772 17076 9824 17128
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 5356 17008 5408 17060
rect 6736 16940 6788 16992
rect 7012 16983 7064 16992
rect 7012 16949 7021 16983
rect 7021 16949 7055 16983
rect 7055 16949 7064 16983
rect 7012 16940 7064 16949
rect 9680 17008 9732 17060
rect 12256 17144 12308 17196
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 13452 17187 13504 17196
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 17776 17212 17828 17264
rect 14464 17076 14516 17128
rect 12164 17008 12216 17060
rect 13636 17008 13688 17060
rect 13728 17008 13780 17060
rect 16120 17076 16172 17128
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 19984 17212 20036 17264
rect 23388 17255 23440 17264
rect 23388 17221 23422 17255
rect 23422 17221 23440 17255
rect 23388 17212 23440 17221
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 21364 17144 21416 17196
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 19524 17076 19576 17128
rect 24768 17144 24820 17196
rect 25504 17187 25556 17196
rect 25504 17153 25513 17187
rect 25513 17153 25547 17187
rect 25547 17153 25556 17187
rect 25504 17144 25556 17153
rect 25596 17144 25648 17196
rect 9404 16940 9456 16992
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10968 16983 11020 16992
rect 10968 16949 10977 16983
rect 10977 16949 11011 16983
rect 11011 16949 11020 16983
rect 10968 16940 11020 16949
rect 11796 16940 11848 16992
rect 12624 16940 12676 16992
rect 15016 16940 15068 16992
rect 16028 16940 16080 16992
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 17776 16940 17828 16949
rect 19984 17008 20036 17060
rect 21456 17008 21508 17060
rect 19800 16940 19852 16992
rect 19892 16940 19944 16992
rect 20720 16940 20772 16992
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 26240 17280 26292 17332
rect 26332 17280 26384 17332
rect 26608 17323 26660 17332
rect 26608 17289 26617 17323
rect 26617 17289 26651 17323
rect 26651 17289 26660 17323
rect 26608 17280 26660 17289
rect 30380 17212 30432 17264
rect 26240 17187 26292 17196
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 28264 17144 28316 17196
rect 30012 17144 30064 17196
rect 24952 17008 25004 17060
rect 22100 16940 22152 16992
rect 25688 17008 25740 17060
rect 27252 17076 27304 17128
rect 28816 17119 28868 17128
rect 28816 17085 28825 17119
rect 28825 17085 28859 17119
rect 28859 17085 28868 17119
rect 28816 17076 28868 17085
rect 29092 17076 29144 17128
rect 30288 17119 30340 17128
rect 30288 17085 30297 17119
rect 30297 17085 30331 17119
rect 30331 17085 30340 17119
rect 30288 17076 30340 17085
rect 25504 16940 25556 16992
rect 26148 16940 26200 16992
rect 27620 16940 27672 16992
rect 28908 16940 28960 16992
rect 30472 16940 30524 16992
rect 4871 16838 4923 16890
rect 4935 16838 4987 16890
rect 4999 16838 5051 16890
rect 5063 16838 5115 16890
rect 5127 16838 5179 16890
rect 12713 16838 12765 16890
rect 12777 16838 12829 16890
rect 12841 16838 12893 16890
rect 12905 16838 12957 16890
rect 12969 16838 13021 16890
rect 20555 16838 20607 16890
rect 20619 16838 20671 16890
rect 20683 16838 20735 16890
rect 20747 16838 20799 16890
rect 20811 16838 20863 16890
rect 28397 16838 28449 16890
rect 28461 16838 28513 16890
rect 28525 16838 28577 16890
rect 28589 16838 28641 16890
rect 28653 16838 28705 16890
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 2688 16600 2740 16652
rect 3056 16643 3108 16652
rect 3056 16609 3065 16643
rect 3065 16609 3099 16643
rect 3099 16609 3108 16643
rect 3056 16600 3108 16609
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 3148 16600 3200 16609
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 4160 16736 4212 16788
rect 8116 16736 8168 16788
rect 10048 16736 10100 16788
rect 12440 16736 12492 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 14740 16736 14792 16788
rect 15752 16736 15804 16788
rect 16028 16736 16080 16788
rect 7196 16668 7248 16720
rect 3240 16600 3292 16609
rect 2320 16507 2372 16516
rect 2320 16473 2329 16507
rect 2329 16473 2363 16507
rect 2363 16473 2372 16507
rect 2320 16464 2372 16473
rect 2872 16396 2924 16448
rect 3608 16532 3660 16584
rect 9312 16668 9364 16720
rect 9404 16668 9456 16720
rect 8208 16600 8260 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10232 16600 10284 16652
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 12624 16668 12676 16720
rect 13452 16668 13504 16720
rect 14832 16668 14884 16720
rect 11428 16600 11480 16652
rect 4252 16507 4304 16516
rect 4252 16473 4286 16507
rect 4286 16473 4304 16507
rect 4252 16464 4304 16473
rect 4344 16396 4396 16448
rect 5264 16464 5316 16516
rect 7288 16464 7340 16516
rect 9956 16532 10008 16584
rect 10416 16464 10468 16516
rect 10784 16575 10836 16584
rect 10784 16541 10793 16575
rect 10793 16541 10827 16575
rect 10827 16541 10836 16575
rect 10784 16532 10836 16541
rect 11612 16532 11664 16584
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 13360 16600 13412 16652
rect 14372 16600 14424 16652
rect 15108 16600 15160 16652
rect 20904 16736 20956 16788
rect 21088 16668 21140 16720
rect 12256 16532 12308 16584
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 13452 16532 13504 16584
rect 14832 16575 14884 16584
rect 14832 16541 14841 16575
rect 14841 16541 14875 16575
rect 14875 16541 14884 16575
rect 14832 16532 14884 16541
rect 15660 16532 15712 16584
rect 19432 16600 19484 16652
rect 21272 16600 21324 16652
rect 21916 16600 21968 16652
rect 23112 16736 23164 16788
rect 24308 16736 24360 16788
rect 25228 16736 25280 16788
rect 26516 16736 26568 16788
rect 29092 16736 29144 16788
rect 31116 16779 31168 16788
rect 31116 16745 31125 16779
rect 31125 16745 31159 16779
rect 31159 16745 31168 16779
rect 31116 16736 31168 16745
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 19708 16532 19760 16584
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 15936 16464 15988 16516
rect 19432 16464 19484 16516
rect 19800 16507 19852 16516
rect 19800 16473 19809 16507
rect 19809 16473 19843 16507
rect 19843 16473 19852 16507
rect 19800 16464 19852 16473
rect 7012 16396 7064 16448
rect 9680 16396 9732 16448
rect 11428 16396 11480 16448
rect 13084 16396 13136 16448
rect 17500 16439 17552 16448
rect 17500 16405 17509 16439
rect 17509 16405 17543 16439
rect 17543 16405 17552 16439
rect 17500 16396 17552 16405
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 20996 16507 21048 16516
rect 20996 16473 21005 16507
rect 21005 16473 21039 16507
rect 21039 16473 21048 16507
rect 20996 16464 21048 16473
rect 21180 16507 21232 16516
rect 21180 16473 21189 16507
rect 21189 16473 21223 16507
rect 21223 16473 21232 16507
rect 21180 16464 21232 16473
rect 22100 16532 22152 16584
rect 28264 16711 28316 16720
rect 28264 16677 28273 16711
rect 28273 16677 28307 16711
rect 28307 16677 28316 16711
rect 28264 16668 28316 16677
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 25136 16600 25188 16652
rect 24124 16532 24176 16584
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 26056 16600 26108 16652
rect 26424 16600 26476 16652
rect 20076 16396 20128 16448
rect 22284 16396 22336 16448
rect 25228 16464 25280 16516
rect 26056 16507 26108 16516
rect 26056 16473 26065 16507
rect 26065 16473 26099 16507
rect 26099 16473 26108 16507
rect 26056 16464 26108 16473
rect 28172 16464 28224 16516
rect 28632 16507 28684 16516
rect 28632 16473 28641 16507
rect 28641 16473 28675 16507
rect 28675 16473 28684 16507
rect 28632 16464 28684 16473
rect 23940 16439 23992 16448
rect 23940 16405 23949 16439
rect 23949 16405 23983 16439
rect 23983 16405 23992 16439
rect 23940 16396 23992 16405
rect 24400 16396 24452 16448
rect 26240 16396 26292 16448
rect 29828 16532 29880 16584
rect 31852 16575 31904 16584
rect 31852 16541 31861 16575
rect 31861 16541 31895 16575
rect 31895 16541 31904 16575
rect 31852 16532 31904 16541
rect 31668 16439 31720 16448
rect 31668 16405 31677 16439
rect 31677 16405 31711 16439
rect 31711 16405 31720 16439
rect 31668 16396 31720 16405
rect 8792 16294 8844 16346
rect 8856 16294 8908 16346
rect 8920 16294 8972 16346
rect 8984 16294 9036 16346
rect 9048 16294 9100 16346
rect 16634 16294 16686 16346
rect 16698 16294 16750 16346
rect 16762 16294 16814 16346
rect 16826 16294 16878 16346
rect 16890 16294 16942 16346
rect 24476 16294 24528 16346
rect 24540 16294 24592 16346
rect 24604 16294 24656 16346
rect 24668 16294 24720 16346
rect 24732 16294 24784 16346
rect 32318 16294 32370 16346
rect 32382 16294 32434 16346
rect 32446 16294 32498 16346
rect 32510 16294 32562 16346
rect 32574 16294 32626 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 2320 16124 2372 16176
rect 2044 16056 2096 16108
rect 3792 16099 3844 16108
rect 3792 16065 3801 16099
rect 3801 16065 3835 16099
rect 3835 16065 3844 16099
rect 3792 16056 3844 16065
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 5080 16235 5132 16244
rect 5080 16201 5089 16235
rect 5089 16201 5123 16235
rect 5123 16201 5132 16235
rect 5080 16192 5132 16201
rect 4068 16124 4120 16176
rect 8392 16192 8444 16244
rect 10968 16192 11020 16244
rect 12532 16192 12584 16244
rect 15660 16192 15712 16244
rect 4068 15988 4120 16040
rect 6092 16056 6144 16108
rect 7104 16124 7156 16176
rect 9588 16167 9640 16176
rect 9588 16133 9597 16167
rect 9597 16133 9631 16167
rect 9631 16133 9640 16167
rect 9588 16124 9640 16133
rect 10324 16124 10376 16176
rect 13360 16124 13412 16176
rect 14648 16167 14700 16176
rect 14648 16133 14657 16167
rect 14657 16133 14691 16167
rect 14691 16133 14700 16167
rect 14648 16124 14700 16133
rect 16120 16124 16172 16176
rect 18420 16167 18472 16176
rect 18420 16133 18429 16167
rect 18429 16133 18463 16167
rect 18463 16133 18472 16167
rect 18420 16124 18472 16133
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 3608 15920 3660 15972
rect 5080 15920 5132 15972
rect 5264 15963 5316 15972
rect 5264 15929 5273 15963
rect 5273 15929 5307 15963
rect 5307 15929 5316 15963
rect 5264 15920 5316 15929
rect 9220 16056 9272 16108
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 11980 16099 12032 16108
rect 8300 15988 8352 16040
rect 8392 15988 8444 16040
rect 8484 15920 8536 15972
rect 10600 15963 10652 15972
rect 10600 15929 10609 15963
rect 10609 15929 10643 15963
rect 10643 15929 10652 15963
rect 10600 15920 10652 15929
rect 11520 15988 11572 16040
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 13084 16056 13136 16108
rect 13452 16056 13504 16108
rect 15476 16056 15528 16108
rect 12072 15988 12124 16040
rect 12164 15988 12216 16040
rect 15844 15988 15896 16040
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 17776 16056 17828 16108
rect 19616 16192 19668 16244
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 19984 16192 20036 16244
rect 20168 16192 20220 16244
rect 24032 16192 24084 16244
rect 25596 16192 25648 16244
rect 28632 16192 28684 16244
rect 29736 16235 29788 16244
rect 29736 16201 29745 16235
rect 29745 16201 29779 16235
rect 29779 16201 29788 16235
rect 29736 16192 29788 16201
rect 31944 16192 31996 16244
rect 20076 16056 20128 16108
rect 19892 15988 19944 16040
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 20904 16056 20956 16065
rect 23204 16124 23256 16176
rect 24124 16124 24176 16176
rect 25044 16056 25096 16108
rect 25412 16056 25464 16108
rect 26608 16124 26660 16176
rect 27620 16124 27672 16176
rect 21732 15988 21784 16040
rect 12992 15920 13044 15972
rect 18880 15920 18932 15972
rect 7472 15852 7524 15904
rect 8116 15852 8168 15904
rect 9220 15852 9272 15904
rect 10508 15852 10560 15904
rect 10692 15852 10744 15904
rect 11336 15852 11388 15904
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 13176 15852 13228 15904
rect 16488 15852 16540 15904
rect 19248 15852 19300 15904
rect 19524 15920 19576 15972
rect 20996 15852 21048 15904
rect 21088 15852 21140 15904
rect 23664 15920 23716 15972
rect 24308 15920 24360 15972
rect 25872 16031 25924 16040
rect 25872 15997 25881 16031
rect 25881 15997 25915 16031
rect 25915 15997 25924 16031
rect 25872 15988 25924 15997
rect 26332 16099 26384 16108
rect 26332 16065 26341 16099
rect 26341 16065 26375 16099
rect 26375 16065 26384 16099
rect 26332 16056 26384 16065
rect 28172 16056 28224 16108
rect 28908 16056 28960 16108
rect 30380 16124 30432 16176
rect 31024 16056 31076 16108
rect 25136 15920 25188 15972
rect 29276 15988 29328 16040
rect 31116 16031 31168 16040
rect 31116 15997 31125 16031
rect 31125 15997 31159 16031
rect 31159 15997 31168 16031
rect 31116 15988 31168 15997
rect 22744 15852 22796 15904
rect 22928 15852 22980 15904
rect 24952 15852 25004 15904
rect 28172 15852 28224 15904
rect 4871 15750 4923 15802
rect 4935 15750 4987 15802
rect 4999 15750 5051 15802
rect 5063 15750 5115 15802
rect 5127 15750 5179 15802
rect 12713 15750 12765 15802
rect 12777 15750 12829 15802
rect 12841 15750 12893 15802
rect 12905 15750 12957 15802
rect 12969 15750 13021 15802
rect 20555 15750 20607 15802
rect 20619 15750 20671 15802
rect 20683 15750 20735 15802
rect 20747 15750 20799 15802
rect 20811 15750 20863 15802
rect 28397 15750 28449 15802
rect 28461 15750 28513 15802
rect 28525 15750 28577 15802
rect 28589 15750 28641 15802
rect 28653 15750 28705 15802
rect 6092 15691 6144 15700
rect 6092 15657 6101 15691
rect 6101 15657 6135 15691
rect 6135 15657 6144 15691
rect 6092 15648 6144 15657
rect 8392 15648 8444 15700
rect 8576 15648 8628 15700
rect 11244 15648 11296 15700
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 2872 15580 2924 15632
rect 3608 15580 3660 15632
rect 10692 15580 10744 15632
rect 11612 15580 11664 15632
rect 14372 15623 14424 15632
rect 14372 15589 14381 15623
rect 14381 15589 14415 15623
rect 14415 15589 14424 15623
rect 14372 15580 14424 15589
rect 15108 15691 15160 15700
rect 15108 15657 15117 15691
rect 15117 15657 15151 15691
rect 15151 15657 15160 15691
rect 15108 15648 15160 15657
rect 16488 15648 16540 15700
rect 17684 15648 17736 15700
rect 18512 15648 18564 15700
rect 19616 15648 19668 15700
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21364 15648 21416 15700
rect 21824 15691 21876 15700
rect 21824 15657 21833 15691
rect 21833 15657 21867 15691
rect 21867 15657 21876 15691
rect 21824 15648 21876 15657
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 25044 15691 25096 15700
rect 25044 15657 25053 15691
rect 25053 15657 25087 15691
rect 25087 15657 25096 15691
rect 25044 15648 25096 15657
rect 25320 15648 25372 15700
rect 4068 15512 4120 15564
rect 7472 15555 7524 15564
rect 7472 15521 7481 15555
rect 7481 15521 7515 15555
rect 7515 15521 7524 15555
rect 7472 15512 7524 15521
rect 11244 15512 11296 15564
rect 11520 15512 11572 15564
rect 12624 15512 12676 15564
rect 3240 15444 3292 15496
rect 3792 15444 3844 15496
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 10140 15444 10192 15496
rect 3516 15376 3568 15428
rect 8392 15376 8444 15428
rect 8576 15376 8628 15428
rect 11888 15444 11940 15496
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 12256 15444 12308 15496
rect 13636 15444 13688 15496
rect 15200 15444 15252 15496
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 18696 15512 18748 15564
rect 21732 15580 21784 15632
rect 27436 15648 27488 15700
rect 28540 15648 28592 15700
rect 19156 15512 19208 15564
rect 11520 15419 11572 15428
rect 11520 15385 11529 15419
rect 11529 15385 11563 15419
rect 11563 15385 11572 15419
rect 11520 15376 11572 15385
rect 13360 15419 13412 15428
rect 13360 15385 13369 15419
rect 13369 15385 13403 15419
rect 13403 15385 13412 15419
rect 13360 15376 13412 15385
rect 13912 15376 13964 15428
rect 14464 15376 14516 15428
rect 2136 15308 2188 15360
rect 3608 15308 3660 15360
rect 10600 15308 10652 15360
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 15476 15308 15528 15360
rect 16488 15308 16540 15360
rect 17316 15308 17368 15360
rect 17776 15351 17828 15360
rect 17776 15317 17803 15351
rect 17803 15317 17828 15351
rect 17776 15308 17828 15317
rect 18420 15376 18472 15428
rect 19248 15444 19300 15496
rect 20168 15512 20220 15564
rect 19616 15444 19668 15496
rect 20904 15512 20956 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 20444 15444 20496 15496
rect 20996 15487 21048 15496
rect 20996 15453 21005 15487
rect 21005 15453 21039 15487
rect 21039 15453 21048 15487
rect 22928 15512 22980 15564
rect 20996 15444 21048 15453
rect 21640 15444 21692 15496
rect 22284 15444 22336 15496
rect 23204 15512 23256 15564
rect 23664 15555 23716 15564
rect 23664 15521 23674 15555
rect 23674 15521 23708 15555
rect 23708 15521 23716 15555
rect 23664 15512 23716 15521
rect 25780 15580 25832 15632
rect 26792 15580 26844 15632
rect 29276 15648 29328 15700
rect 31024 15691 31076 15700
rect 31024 15657 31033 15691
rect 31033 15657 31067 15691
rect 31067 15657 31076 15691
rect 31024 15648 31076 15657
rect 23940 15512 23992 15564
rect 30196 15512 30248 15564
rect 30380 15580 30432 15632
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 23756 15444 23808 15496
rect 20812 15376 20864 15428
rect 21732 15419 21784 15428
rect 21732 15385 21741 15419
rect 21741 15385 21775 15419
rect 21775 15385 21784 15419
rect 21732 15376 21784 15385
rect 18328 15308 18380 15360
rect 18604 15308 18656 15360
rect 19156 15308 19208 15360
rect 20260 15308 20312 15360
rect 20352 15351 20404 15360
rect 20352 15317 20361 15351
rect 20361 15317 20395 15351
rect 20395 15317 20404 15351
rect 20352 15308 20404 15317
rect 22744 15376 22796 15428
rect 24860 15376 24912 15428
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 25320 15487 25372 15496
rect 25320 15453 25329 15487
rect 25329 15453 25363 15487
rect 25363 15453 25372 15487
rect 25320 15444 25372 15453
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 25688 15444 25740 15496
rect 26056 15487 26108 15496
rect 26056 15453 26065 15487
rect 26065 15453 26099 15487
rect 26099 15453 26108 15487
rect 26056 15444 26108 15453
rect 29000 15444 29052 15496
rect 30012 15444 30064 15496
rect 30104 15376 30156 15428
rect 24308 15308 24360 15360
rect 27436 15308 27488 15360
rect 27712 15308 27764 15360
rect 28540 15308 28592 15360
rect 30380 15308 30432 15360
rect 31668 15308 31720 15360
rect 8792 15206 8844 15258
rect 8856 15206 8908 15258
rect 8920 15206 8972 15258
rect 8984 15206 9036 15258
rect 9048 15206 9100 15258
rect 16634 15206 16686 15258
rect 16698 15206 16750 15258
rect 16762 15206 16814 15258
rect 16826 15206 16878 15258
rect 16890 15206 16942 15258
rect 24476 15206 24528 15258
rect 24540 15206 24592 15258
rect 24604 15206 24656 15258
rect 24668 15206 24720 15258
rect 24732 15206 24784 15258
rect 32318 15206 32370 15258
rect 32382 15206 32434 15258
rect 32446 15206 32498 15258
rect 32510 15206 32562 15258
rect 32574 15206 32626 15258
rect 8576 15104 8628 15156
rect 16120 15147 16172 15156
rect 16120 15113 16129 15147
rect 16129 15113 16163 15147
rect 16163 15113 16172 15147
rect 16120 15104 16172 15113
rect 9956 15036 10008 15088
rect 11428 15036 11480 15088
rect 11980 15036 12032 15088
rect 3056 14968 3108 15020
rect 3976 14968 4028 15020
rect 7104 14968 7156 15020
rect 8484 14968 8536 15020
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 11704 14968 11756 15020
rect 12440 14968 12492 15020
rect 13544 14968 13596 15020
rect 13636 15011 13688 15020
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 13912 15011 13964 15020
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 14372 14968 14424 15020
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 17776 15104 17828 15156
rect 18512 15147 18564 15156
rect 18512 15113 18521 15147
rect 18521 15113 18555 15147
rect 18555 15113 18564 15147
rect 18512 15104 18564 15113
rect 22192 15104 22244 15156
rect 16488 14968 16540 15020
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 20812 15079 20864 15088
rect 20812 15045 20821 15079
rect 20821 15045 20855 15079
rect 20855 15045 20864 15079
rect 20812 15036 20864 15045
rect 21456 15036 21508 15088
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 2596 14900 2648 14909
rect 6092 14900 6144 14952
rect 6644 14900 6696 14952
rect 13360 14900 13412 14952
rect 13728 14900 13780 14952
rect 14096 14943 14148 14952
rect 14096 14909 14105 14943
rect 14105 14909 14139 14943
rect 14139 14909 14148 14943
rect 14096 14900 14148 14909
rect 17776 15011 17828 15020
rect 17776 14977 17785 15011
rect 17785 14977 17819 15011
rect 17819 14977 17828 15011
rect 17776 14968 17828 14977
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 19248 14968 19300 15020
rect 20168 14968 20220 15020
rect 20444 14968 20496 15020
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 23572 15036 23624 15088
rect 24216 15104 24268 15156
rect 24952 15104 25004 15156
rect 26240 15104 26292 15156
rect 28724 15104 28776 15156
rect 29736 15104 29788 15156
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23296 14968 23348 15020
rect 25136 15036 25188 15088
rect 27436 15036 27488 15088
rect 28080 15036 28132 15088
rect 28264 15036 28316 15088
rect 30012 15036 30064 15088
rect 31116 15036 31168 15088
rect 24860 14968 24912 15020
rect 25780 15011 25832 15020
rect 25780 14977 25789 15011
rect 25789 14977 25823 15011
rect 25823 14977 25832 15011
rect 25780 14968 25832 14977
rect 25964 14968 26016 15020
rect 26332 14968 26384 15020
rect 26516 14968 26568 15020
rect 5632 14832 5684 14884
rect 6920 14832 6972 14884
rect 10140 14875 10192 14884
rect 10140 14841 10149 14875
rect 10149 14841 10183 14875
rect 10183 14841 10192 14875
rect 10140 14832 10192 14841
rect 11888 14832 11940 14884
rect 14648 14832 14700 14884
rect 4528 14764 4580 14816
rect 8116 14764 8168 14816
rect 9312 14764 9364 14816
rect 9588 14807 9640 14816
rect 9588 14773 9597 14807
rect 9597 14773 9631 14807
rect 9631 14773 9640 14807
rect 9588 14764 9640 14773
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 10692 14807 10744 14816
rect 10692 14773 10701 14807
rect 10701 14773 10735 14807
rect 10735 14773 10744 14807
rect 10692 14764 10744 14773
rect 13636 14764 13688 14816
rect 18604 14900 18656 14952
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 18788 14943 18840 14952
rect 18788 14909 18797 14943
rect 18797 14909 18831 14943
rect 18831 14909 18840 14943
rect 18788 14900 18840 14909
rect 15752 14832 15804 14884
rect 17040 14832 17092 14884
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 19156 14900 19208 14952
rect 19708 14943 19760 14952
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 16304 14807 16356 14816
rect 16304 14773 16313 14807
rect 16313 14773 16347 14807
rect 16347 14773 16356 14807
rect 16304 14764 16356 14773
rect 16948 14764 17000 14816
rect 17132 14764 17184 14816
rect 19984 14832 20036 14884
rect 21640 14900 21692 14952
rect 20260 14764 20312 14816
rect 22468 14764 22520 14816
rect 25872 14900 25924 14952
rect 28908 14900 28960 14952
rect 29368 15011 29420 15020
rect 29368 14977 29377 15011
rect 29377 14977 29411 15011
rect 29411 14977 29420 15011
rect 29368 14968 29420 14977
rect 30472 14968 30524 15020
rect 31392 15011 31444 15020
rect 31392 14977 31410 15011
rect 31410 14977 31444 15011
rect 31392 14968 31444 14977
rect 29552 14900 29604 14952
rect 23940 14764 23992 14816
rect 25320 14764 25372 14816
rect 25688 14764 25740 14816
rect 26608 14764 26660 14816
rect 27528 14764 27580 14816
rect 28172 14807 28224 14816
rect 28172 14773 28181 14807
rect 28181 14773 28215 14807
rect 28215 14773 28224 14807
rect 28172 14764 28224 14773
rect 29644 14807 29696 14816
rect 29644 14773 29653 14807
rect 29653 14773 29687 14807
rect 29687 14773 29696 14807
rect 29644 14764 29696 14773
rect 29828 14807 29880 14816
rect 29828 14773 29837 14807
rect 29837 14773 29871 14807
rect 29871 14773 29880 14807
rect 29828 14764 29880 14773
rect 4871 14662 4923 14714
rect 4935 14662 4987 14714
rect 4999 14662 5051 14714
rect 5063 14662 5115 14714
rect 5127 14662 5179 14714
rect 12713 14662 12765 14714
rect 12777 14662 12829 14714
rect 12841 14662 12893 14714
rect 12905 14662 12957 14714
rect 12969 14662 13021 14714
rect 20555 14662 20607 14714
rect 20619 14662 20671 14714
rect 20683 14662 20735 14714
rect 20747 14662 20799 14714
rect 20811 14662 20863 14714
rect 28397 14662 28449 14714
rect 28461 14662 28513 14714
rect 28525 14662 28577 14714
rect 28589 14662 28641 14714
rect 28653 14662 28705 14714
rect 3148 14560 3200 14612
rect 8300 14560 8352 14612
rect 8392 14603 8444 14612
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 6368 14492 6420 14544
rect 7656 14424 7708 14476
rect 8300 14424 8352 14476
rect 9772 14492 9824 14544
rect 10784 14560 10836 14612
rect 12072 14560 12124 14612
rect 12716 14603 12768 14612
rect 12716 14569 12725 14603
rect 12725 14569 12759 14603
rect 12759 14569 12768 14603
rect 12716 14560 12768 14569
rect 2412 14356 2464 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 7104 14356 7156 14408
rect 8116 14356 8168 14408
rect 3516 14288 3568 14340
rect 7656 14288 7708 14340
rect 9588 14356 9640 14408
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 13452 14560 13504 14612
rect 14188 14424 14240 14476
rect 14648 14560 14700 14612
rect 11428 14288 11480 14340
rect 3056 14220 3108 14272
rect 3424 14220 3476 14272
rect 3700 14220 3752 14272
rect 4436 14220 4488 14272
rect 6736 14220 6788 14272
rect 9680 14220 9732 14272
rect 11612 14331 11664 14340
rect 11612 14297 11630 14331
rect 11630 14297 11664 14331
rect 11612 14288 11664 14297
rect 12716 14331 12768 14340
rect 12716 14297 12725 14331
rect 12725 14297 12759 14331
rect 12759 14297 12768 14331
rect 12716 14288 12768 14297
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 13636 14288 13688 14340
rect 14372 14356 14424 14408
rect 15384 14356 15436 14408
rect 16304 14356 16356 14408
rect 21732 14560 21784 14612
rect 21824 14560 21876 14612
rect 23296 14560 23348 14612
rect 24308 14560 24360 14612
rect 25136 14603 25188 14612
rect 25136 14569 25145 14603
rect 25145 14569 25179 14603
rect 25179 14569 25188 14603
rect 25136 14560 25188 14569
rect 25228 14560 25280 14612
rect 22192 14467 22244 14476
rect 22192 14433 22201 14467
rect 22201 14433 22235 14467
rect 22235 14433 22244 14467
rect 22192 14424 22244 14433
rect 22560 14424 22612 14476
rect 23112 14424 23164 14476
rect 19800 14399 19852 14408
rect 19800 14365 19809 14399
rect 19809 14365 19843 14399
rect 19843 14365 19852 14399
rect 19800 14356 19852 14365
rect 20352 14356 20404 14408
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 18788 14288 18840 14340
rect 12440 14220 12492 14272
rect 13820 14220 13872 14272
rect 15292 14220 15344 14272
rect 15936 14220 15988 14272
rect 17408 14220 17460 14272
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 18972 14220 19024 14272
rect 21824 14220 21876 14272
rect 24400 14356 24452 14408
rect 24952 14399 25004 14408
rect 24952 14365 24961 14399
rect 24961 14365 24995 14399
rect 24995 14365 25004 14399
rect 24952 14356 25004 14365
rect 25136 14356 25188 14408
rect 25780 14424 25832 14476
rect 25872 14399 25924 14408
rect 25872 14365 25881 14399
rect 25881 14365 25915 14399
rect 25915 14365 25924 14399
rect 25872 14356 25924 14365
rect 26240 14560 26292 14612
rect 28172 14560 28224 14612
rect 26332 14492 26384 14544
rect 26608 14424 26660 14476
rect 27712 14424 27764 14476
rect 28816 14424 28868 14476
rect 31116 14560 31168 14612
rect 26240 14356 26292 14408
rect 27436 14356 27488 14408
rect 28908 14399 28960 14408
rect 28908 14365 28917 14399
rect 28917 14365 28951 14399
rect 28951 14365 28960 14399
rect 28908 14356 28960 14365
rect 29828 14356 29880 14408
rect 25412 14288 25464 14340
rect 25964 14331 26016 14340
rect 25964 14297 25973 14331
rect 25973 14297 26007 14331
rect 26007 14297 26016 14331
rect 25964 14288 26016 14297
rect 28816 14331 28868 14340
rect 28816 14297 28825 14331
rect 28825 14297 28859 14331
rect 28859 14297 28868 14331
rect 28816 14288 28868 14297
rect 23848 14220 23900 14272
rect 24216 14220 24268 14272
rect 24952 14220 25004 14272
rect 25320 14220 25372 14272
rect 26148 14220 26200 14272
rect 26240 14263 26292 14272
rect 26240 14229 26249 14263
rect 26249 14229 26283 14263
rect 26283 14229 26292 14263
rect 26240 14220 26292 14229
rect 28080 14263 28132 14272
rect 28080 14229 28089 14263
rect 28089 14229 28123 14263
rect 28123 14229 28132 14263
rect 28080 14220 28132 14229
rect 28724 14220 28776 14272
rect 30104 14288 30156 14340
rect 29736 14220 29788 14272
rect 8792 14118 8844 14170
rect 8856 14118 8908 14170
rect 8920 14118 8972 14170
rect 8984 14118 9036 14170
rect 9048 14118 9100 14170
rect 16634 14118 16686 14170
rect 16698 14118 16750 14170
rect 16762 14118 16814 14170
rect 16826 14118 16878 14170
rect 16890 14118 16942 14170
rect 24476 14118 24528 14170
rect 24540 14118 24592 14170
rect 24604 14118 24656 14170
rect 24668 14118 24720 14170
rect 24732 14118 24784 14170
rect 32318 14118 32370 14170
rect 32382 14118 32434 14170
rect 32446 14118 32498 14170
rect 32510 14118 32562 14170
rect 32574 14118 32626 14170
rect 3516 14016 3568 14068
rect 9680 14016 9732 14068
rect 10508 14016 10560 14068
rect 11612 14016 11664 14068
rect 12716 14016 12768 14068
rect 3700 13948 3752 14000
rect 5632 13991 5684 14000
rect 5632 13957 5641 13991
rect 5641 13957 5675 13991
rect 5675 13957 5684 13991
rect 5632 13948 5684 13957
rect 6736 13948 6788 14000
rect 7748 13948 7800 14000
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9312 13880 9364 13932
rect 10692 13880 10744 13932
rect 13820 13880 13872 13932
rect 14832 14016 14884 14068
rect 15568 14016 15620 14068
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 23388 14016 23440 14068
rect 26056 14016 26108 14068
rect 15292 13991 15344 14000
rect 15292 13957 15301 13991
rect 15301 13957 15335 13991
rect 15335 13957 15344 13991
rect 15292 13948 15344 13957
rect 16120 13948 16172 14000
rect 31760 14016 31812 14068
rect 28908 13948 28960 14000
rect 30472 13991 30524 14000
rect 30472 13957 30497 13991
rect 30497 13957 30524 13991
rect 30472 13948 30524 13957
rect 15384 13880 15436 13932
rect 15660 13880 15712 13932
rect 17040 13880 17092 13932
rect 17316 13923 17368 13932
rect 17316 13889 17325 13923
rect 17325 13889 17359 13923
rect 17359 13889 17368 13923
rect 17316 13880 17368 13889
rect 21732 13880 21784 13932
rect 22192 13880 22244 13932
rect 4252 13812 4304 13864
rect 4436 13855 4488 13864
rect 4436 13821 4445 13855
rect 4445 13821 4479 13855
rect 4479 13821 4488 13855
rect 4436 13812 4488 13821
rect 2228 13676 2280 13728
rect 2412 13719 2464 13728
rect 2412 13685 2421 13719
rect 2421 13685 2455 13719
rect 2455 13685 2464 13719
rect 2412 13676 2464 13685
rect 5356 13676 5408 13728
rect 13360 13812 13412 13864
rect 13636 13812 13688 13864
rect 15292 13812 15344 13864
rect 18236 13812 18288 13864
rect 20444 13812 20496 13864
rect 21916 13812 21968 13864
rect 22376 13812 22428 13864
rect 23112 13880 23164 13932
rect 22928 13812 22980 13864
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24400 13880 24452 13932
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 25412 13880 25464 13932
rect 26516 13923 26568 13932
rect 26516 13889 26525 13923
rect 26525 13889 26559 13923
rect 26559 13889 26568 13923
rect 26516 13880 26568 13889
rect 27712 13923 27764 13932
rect 27712 13889 27721 13923
rect 27721 13889 27755 13923
rect 27755 13889 27764 13923
rect 27712 13880 27764 13889
rect 27804 13880 27856 13932
rect 29368 13880 29420 13932
rect 29736 13923 29788 13932
rect 29736 13889 29745 13923
rect 29745 13889 29779 13923
rect 29779 13889 29788 13923
rect 29736 13880 29788 13889
rect 24308 13812 24360 13864
rect 6736 13787 6788 13796
rect 6736 13753 6745 13787
rect 6745 13753 6779 13787
rect 6779 13753 6788 13787
rect 6736 13744 6788 13753
rect 17776 13744 17828 13796
rect 25044 13812 25096 13864
rect 25872 13812 25924 13864
rect 26700 13812 26752 13864
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 6552 13676 6604 13685
rect 8116 13719 8168 13728
rect 8116 13685 8125 13719
rect 8125 13685 8159 13719
rect 8159 13685 8168 13719
rect 8116 13676 8168 13685
rect 12624 13676 12676 13728
rect 14740 13676 14792 13728
rect 14924 13676 14976 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 15844 13676 15896 13728
rect 17408 13676 17460 13728
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 22376 13676 22428 13728
rect 22652 13719 22704 13728
rect 22652 13685 22661 13719
rect 22661 13685 22695 13719
rect 22695 13685 22704 13719
rect 22652 13676 22704 13685
rect 24216 13676 24268 13728
rect 26608 13744 26660 13796
rect 29644 13812 29696 13864
rect 31392 13812 31444 13864
rect 25320 13719 25372 13728
rect 25320 13685 25329 13719
rect 25329 13685 25363 13719
rect 25363 13685 25372 13719
rect 25320 13676 25372 13685
rect 25872 13719 25924 13728
rect 25872 13685 25881 13719
rect 25881 13685 25915 13719
rect 25915 13685 25924 13719
rect 25872 13676 25924 13685
rect 29092 13719 29144 13728
rect 29092 13685 29101 13719
rect 29101 13685 29135 13719
rect 29135 13685 29144 13719
rect 29092 13676 29144 13685
rect 30380 13676 30432 13728
rect 4871 13574 4923 13626
rect 4935 13574 4987 13626
rect 4999 13574 5051 13626
rect 5063 13574 5115 13626
rect 5127 13574 5179 13626
rect 12713 13574 12765 13626
rect 12777 13574 12829 13626
rect 12841 13574 12893 13626
rect 12905 13574 12957 13626
rect 12969 13574 13021 13626
rect 20555 13574 20607 13626
rect 20619 13574 20671 13626
rect 20683 13574 20735 13626
rect 20747 13574 20799 13626
rect 20811 13574 20863 13626
rect 28397 13574 28449 13626
rect 28461 13574 28513 13626
rect 28525 13574 28577 13626
rect 28589 13574 28641 13626
rect 28653 13574 28705 13626
rect 3056 13472 3108 13524
rect 5908 13472 5960 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 8116 13472 8168 13524
rect 2136 13268 2188 13320
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 2412 13200 2464 13252
rect 3332 13200 3384 13252
rect 4252 13336 4304 13388
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 10140 13472 10192 13524
rect 10508 13472 10560 13524
rect 12624 13472 12676 13524
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 6736 13268 6788 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 3240 13132 3292 13184
rect 3424 13132 3476 13184
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 5816 13132 5868 13184
rect 6828 13200 6880 13252
rect 9680 13268 9732 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 9404 13200 9456 13252
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 14648 13472 14700 13524
rect 15384 13472 15436 13524
rect 18972 13472 19024 13524
rect 21548 13472 21600 13524
rect 14096 13404 14148 13456
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 15016 13404 15068 13456
rect 15200 13404 15252 13456
rect 15476 13404 15528 13456
rect 19432 13447 19484 13456
rect 19432 13413 19441 13447
rect 19441 13413 19475 13447
rect 19475 13413 19484 13447
rect 19432 13404 19484 13413
rect 19524 13404 19576 13456
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 10784 13243 10836 13252
rect 10784 13209 10793 13243
rect 10793 13209 10827 13243
rect 10827 13209 10836 13243
rect 10784 13200 10836 13209
rect 18420 13336 18472 13388
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 14924 13268 14976 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15568 13268 15620 13320
rect 17500 13268 17552 13320
rect 16120 13200 16172 13252
rect 17776 13200 17828 13252
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 9312 13132 9364 13184
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 12072 13175 12124 13184
rect 12072 13141 12081 13175
rect 12081 13141 12115 13175
rect 12115 13141 12124 13175
rect 12072 13132 12124 13141
rect 13452 13132 13504 13184
rect 13636 13132 13688 13184
rect 14372 13132 14424 13184
rect 15108 13132 15160 13184
rect 19524 13132 19576 13184
rect 22560 13336 22612 13388
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 21548 13268 21600 13320
rect 25964 13515 26016 13524
rect 25964 13481 25973 13515
rect 25973 13481 26007 13515
rect 26007 13481 26016 13515
rect 25964 13472 26016 13481
rect 26332 13472 26384 13524
rect 27804 13515 27856 13524
rect 27804 13481 27813 13515
rect 27813 13481 27847 13515
rect 27847 13481 27856 13515
rect 27804 13472 27856 13481
rect 28264 13472 28316 13524
rect 26148 13404 26200 13456
rect 29000 13404 29052 13456
rect 24308 13336 24360 13388
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 23296 13200 23348 13252
rect 24216 13268 24268 13320
rect 25320 13268 25372 13320
rect 26240 13336 26292 13388
rect 26332 13336 26384 13388
rect 29552 13472 29604 13524
rect 30932 13472 30984 13524
rect 29184 13447 29236 13456
rect 29184 13413 29193 13447
rect 29193 13413 29227 13447
rect 29227 13413 29236 13447
rect 29184 13404 29236 13413
rect 30012 13404 30064 13456
rect 29460 13336 29512 13388
rect 26516 13268 26568 13320
rect 26792 13268 26844 13320
rect 27620 13311 27672 13320
rect 27620 13277 27629 13311
rect 27629 13277 27663 13311
rect 27663 13277 27672 13311
rect 27620 13268 27672 13277
rect 27804 13268 27856 13320
rect 28724 13268 28776 13320
rect 29000 13268 29052 13320
rect 29920 13268 29972 13320
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 24676 13200 24728 13209
rect 25964 13200 26016 13252
rect 26148 13200 26200 13252
rect 26240 13243 26292 13252
rect 26240 13209 26249 13243
rect 26249 13209 26283 13243
rect 26283 13209 26292 13243
rect 26240 13200 26292 13209
rect 22744 13132 22796 13184
rect 23848 13132 23900 13184
rect 27436 13175 27488 13184
rect 27436 13141 27445 13175
rect 27445 13141 27479 13175
rect 27479 13141 27488 13175
rect 27436 13132 27488 13141
rect 27712 13132 27764 13184
rect 27896 13132 27948 13184
rect 29644 13132 29696 13184
rect 8792 13030 8844 13082
rect 8856 13030 8908 13082
rect 8920 13030 8972 13082
rect 8984 13030 9036 13082
rect 9048 13030 9100 13082
rect 16634 13030 16686 13082
rect 16698 13030 16750 13082
rect 16762 13030 16814 13082
rect 16826 13030 16878 13082
rect 16890 13030 16942 13082
rect 24476 13030 24528 13082
rect 24540 13030 24592 13082
rect 24604 13030 24656 13082
rect 24668 13030 24720 13082
rect 24732 13030 24784 13082
rect 32318 13030 32370 13082
rect 32382 13030 32434 13082
rect 32446 13030 32498 13082
rect 32510 13030 32562 13082
rect 32574 13030 32626 13082
rect 2688 12928 2740 12980
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 2872 12792 2924 12844
rect 3976 12928 4028 12980
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 4068 12860 4120 12912
rect 4436 12860 4488 12912
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 3424 12792 3476 12844
rect 3700 12792 3752 12844
rect 6552 12860 6604 12912
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 2872 12656 2924 12708
rect 3148 12656 3200 12708
rect 3240 12656 3292 12708
rect 3700 12588 3752 12640
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 6460 12792 6512 12844
rect 12164 12860 12216 12912
rect 14556 12860 14608 12912
rect 15660 12928 15712 12980
rect 18328 12971 18380 12980
rect 18328 12937 18337 12971
rect 18337 12937 18371 12971
rect 18371 12937 18380 12971
rect 18328 12928 18380 12937
rect 20352 12928 20404 12980
rect 23296 12928 23348 12980
rect 23664 12971 23716 12980
rect 23664 12937 23673 12971
rect 23673 12937 23707 12971
rect 23707 12937 23716 12971
rect 24676 12971 24728 12980
rect 23664 12928 23716 12937
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 24952 12928 25004 12980
rect 25228 12928 25280 12980
rect 7012 12835 7064 12844
rect 7012 12801 7046 12835
rect 7046 12801 7064 12835
rect 7012 12792 7064 12801
rect 9588 12792 9640 12844
rect 9864 12792 9916 12844
rect 11520 12792 11572 12844
rect 13176 12835 13228 12844
rect 13176 12801 13185 12835
rect 13185 12801 13219 12835
rect 13219 12801 13228 12835
rect 13176 12792 13228 12801
rect 13452 12835 13504 12844
rect 13452 12801 13486 12835
rect 13486 12801 13504 12835
rect 13452 12792 13504 12801
rect 13912 12792 13964 12844
rect 15108 12792 15160 12844
rect 16120 12860 16172 12912
rect 18236 12860 18288 12912
rect 19432 12903 19484 12912
rect 19432 12869 19450 12903
rect 19450 12869 19484 12903
rect 19432 12860 19484 12869
rect 20904 12860 20956 12912
rect 16028 12792 16080 12844
rect 21364 12792 21416 12844
rect 22744 12835 22796 12844
rect 22744 12801 22753 12835
rect 22753 12801 22787 12835
rect 22787 12801 22796 12835
rect 22744 12792 22796 12801
rect 23848 12792 23900 12844
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 5724 12724 5776 12776
rect 6552 12724 6604 12776
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 14464 12656 14516 12708
rect 19800 12724 19852 12776
rect 20904 12724 20956 12776
rect 22100 12724 22152 12776
rect 23204 12767 23256 12776
rect 23204 12733 23213 12767
rect 23213 12733 23247 12767
rect 23247 12733 23256 12767
rect 23204 12724 23256 12733
rect 15200 12656 15252 12708
rect 15936 12656 15988 12708
rect 20444 12656 20496 12708
rect 7380 12588 7432 12640
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 10232 12588 10284 12597
rect 13544 12588 13596 12640
rect 19524 12588 19576 12640
rect 22284 12656 22336 12708
rect 22192 12588 22244 12640
rect 22836 12588 22888 12640
rect 23296 12588 23348 12640
rect 25504 12860 25556 12912
rect 26148 12928 26200 12980
rect 27436 12971 27488 12980
rect 27436 12937 27445 12971
rect 27445 12937 27479 12971
rect 27479 12937 27488 12971
rect 27436 12928 27488 12937
rect 29000 12928 29052 12980
rect 29184 12860 29236 12912
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 25596 12724 25648 12776
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 25964 12724 26016 12776
rect 27252 12792 27304 12844
rect 27712 12792 27764 12844
rect 28908 12792 28960 12844
rect 32036 12860 32088 12912
rect 29644 12835 29696 12844
rect 29644 12801 29653 12835
rect 29653 12801 29687 12835
rect 29687 12801 29696 12835
rect 29644 12792 29696 12801
rect 29828 12835 29880 12844
rect 29828 12801 29837 12835
rect 29837 12801 29871 12835
rect 29871 12801 29880 12835
rect 29828 12792 29880 12801
rect 30564 12835 30616 12844
rect 30564 12801 30598 12835
rect 30598 12801 30616 12835
rect 30564 12792 30616 12801
rect 27896 12724 27948 12776
rect 29000 12724 29052 12776
rect 30288 12767 30340 12776
rect 30288 12733 30297 12767
rect 30297 12733 30331 12767
rect 30331 12733 30340 12767
rect 30288 12724 30340 12733
rect 27620 12699 27672 12708
rect 27620 12665 27629 12699
rect 27629 12665 27663 12699
rect 27663 12665 27672 12699
rect 27620 12656 27672 12665
rect 27988 12656 28040 12708
rect 29920 12588 29972 12640
rect 4871 12486 4923 12538
rect 4935 12486 4987 12538
rect 4999 12486 5051 12538
rect 5063 12486 5115 12538
rect 5127 12486 5179 12538
rect 12713 12486 12765 12538
rect 12777 12486 12829 12538
rect 12841 12486 12893 12538
rect 12905 12486 12957 12538
rect 12969 12486 13021 12538
rect 20555 12486 20607 12538
rect 20619 12486 20671 12538
rect 20683 12486 20735 12538
rect 20747 12486 20799 12538
rect 20811 12486 20863 12538
rect 28397 12486 28449 12538
rect 28461 12486 28513 12538
rect 28525 12486 28577 12538
rect 28589 12486 28641 12538
rect 28653 12486 28705 12538
rect 3148 12384 3200 12436
rect 5632 12384 5684 12436
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 13544 12427 13596 12436
rect 13544 12393 13553 12427
rect 13553 12393 13587 12427
rect 13587 12393 13596 12427
rect 13544 12384 13596 12393
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 15384 12384 15436 12436
rect 15752 12384 15804 12436
rect 15844 12384 15896 12436
rect 16488 12384 16540 12436
rect 17132 12384 17184 12436
rect 3332 12316 3384 12368
rect 14280 12359 14332 12368
rect 14280 12325 14289 12359
rect 14289 12325 14323 12359
rect 14323 12325 14332 12359
rect 14280 12316 14332 12325
rect 15200 12316 15252 12368
rect 15568 12316 15620 12368
rect 3148 12248 3200 12300
rect 5540 12248 5592 12300
rect 6368 12248 6420 12300
rect 9956 12248 10008 12300
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 3240 12112 3292 12164
rect 9128 12180 9180 12232
rect 11152 12180 11204 12232
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 13636 12180 13688 12232
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15476 12248 15528 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 19432 12180 19484 12232
rect 21548 12427 21600 12436
rect 21548 12393 21557 12427
rect 21557 12393 21591 12427
rect 21591 12393 21600 12427
rect 21548 12384 21600 12393
rect 22836 12384 22888 12436
rect 23204 12427 23256 12436
rect 23204 12393 23213 12427
rect 23213 12393 23247 12427
rect 23247 12393 23256 12427
rect 23204 12384 23256 12393
rect 26240 12384 26292 12436
rect 27712 12427 27764 12436
rect 27712 12393 27721 12427
rect 27721 12393 27755 12427
rect 27755 12393 27764 12427
rect 27712 12384 27764 12393
rect 30564 12384 30616 12436
rect 23296 12316 23348 12368
rect 22284 12248 22336 12300
rect 22560 12291 22612 12300
rect 22560 12257 22569 12291
rect 22569 12257 22603 12291
rect 22603 12257 22612 12291
rect 22560 12248 22612 12257
rect 22744 12180 22796 12232
rect 24676 12316 24728 12368
rect 29828 12316 29880 12368
rect 25504 12248 25556 12300
rect 25964 12291 26016 12300
rect 25964 12257 25973 12291
rect 25973 12257 26007 12291
rect 26007 12257 26016 12291
rect 25964 12248 26016 12257
rect 29460 12248 29512 12300
rect 30012 12291 30064 12300
rect 30012 12257 30021 12291
rect 30021 12257 30055 12291
rect 30055 12257 30064 12291
rect 30012 12248 30064 12257
rect 6368 12155 6420 12164
rect 6368 12121 6395 12155
rect 6395 12121 6420 12155
rect 6368 12112 6420 12121
rect 6644 12112 6696 12164
rect 10416 12155 10468 12164
rect 10416 12121 10450 12155
rect 10450 12121 10468 12155
rect 10416 12112 10468 12121
rect 13452 12112 13504 12164
rect 15200 12112 15252 12164
rect 15292 12155 15344 12164
rect 15292 12121 15301 12155
rect 15301 12121 15335 12155
rect 15335 12121 15344 12155
rect 15292 12112 15344 12121
rect 17040 12112 17092 12164
rect 12440 12044 12492 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 13912 12044 13964 12096
rect 15476 12087 15528 12096
rect 15476 12053 15511 12087
rect 15511 12053 15528 12087
rect 15476 12044 15528 12053
rect 15844 12044 15896 12096
rect 17776 12044 17828 12096
rect 18604 12112 18656 12164
rect 22100 12112 22152 12164
rect 23664 12112 23716 12164
rect 19156 12044 19208 12096
rect 22652 12044 22704 12096
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 25780 12223 25832 12232
rect 25780 12189 25789 12223
rect 25789 12189 25823 12223
rect 25823 12189 25832 12223
rect 25780 12180 25832 12189
rect 25688 12112 25740 12164
rect 26056 12180 26108 12232
rect 29092 12223 29144 12232
rect 29092 12189 29101 12223
rect 29101 12189 29135 12223
rect 29135 12189 29144 12223
rect 29092 12180 29144 12189
rect 29644 12180 29696 12232
rect 25320 12044 25372 12096
rect 28080 12087 28132 12096
rect 28080 12053 28089 12087
rect 28089 12053 28123 12087
rect 28123 12053 28132 12087
rect 28080 12044 28132 12053
rect 28172 12087 28224 12096
rect 28172 12053 28181 12087
rect 28181 12053 28215 12087
rect 28215 12053 28224 12087
rect 28172 12044 28224 12053
rect 29276 12112 29328 12164
rect 30196 12223 30248 12232
rect 30196 12189 30205 12223
rect 30205 12189 30239 12223
rect 30239 12189 30248 12223
rect 30196 12180 30248 12189
rect 30748 12180 30800 12232
rect 30380 12112 30432 12164
rect 29000 12087 29052 12096
rect 29000 12053 29015 12087
rect 29015 12053 29049 12087
rect 29049 12053 29052 12087
rect 29000 12044 29052 12053
rect 29736 12087 29788 12096
rect 29736 12053 29745 12087
rect 29745 12053 29779 12087
rect 29779 12053 29788 12087
rect 29736 12044 29788 12053
rect 8792 11942 8844 11994
rect 8856 11942 8908 11994
rect 8920 11942 8972 11994
rect 8984 11942 9036 11994
rect 9048 11942 9100 11994
rect 16634 11942 16686 11994
rect 16698 11942 16750 11994
rect 16762 11942 16814 11994
rect 16826 11942 16878 11994
rect 16890 11942 16942 11994
rect 24476 11942 24528 11994
rect 24540 11942 24592 11994
rect 24604 11942 24656 11994
rect 24668 11942 24720 11994
rect 24732 11942 24784 11994
rect 32318 11942 32370 11994
rect 32382 11942 32434 11994
rect 32446 11942 32498 11994
rect 32510 11942 32562 11994
rect 32574 11942 32626 11994
rect 2964 11840 3016 11892
rect 4068 11840 4120 11892
rect 14832 11840 14884 11892
rect 15476 11840 15528 11892
rect 2872 11772 2924 11824
rect 7748 11772 7800 11824
rect 12532 11772 12584 11824
rect 14648 11815 14700 11824
rect 14648 11781 14657 11815
rect 14657 11781 14691 11815
rect 14691 11781 14700 11815
rect 14648 11772 14700 11781
rect 15200 11772 15252 11824
rect 15844 11772 15896 11824
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 3608 11704 3660 11756
rect 4712 11704 4764 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 7380 11704 7432 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 14096 11704 14148 11756
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 15568 11704 15620 11756
rect 25780 11840 25832 11892
rect 28172 11883 28224 11892
rect 28172 11849 28181 11883
rect 28181 11849 28215 11883
rect 28215 11849 28224 11883
rect 28172 11840 28224 11849
rect 29368 11883 29420 11892
rect 29368 11849 29377 11883
rect 29377 11849 29411 11883
rect 29411 11849 29420 11883
rect 29368 11840 29420 11849
rect 30196 11840 30248 11892
rect 17868 11772 17920 11824
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 17224 11704 17276 11756
rect 17776 11747 17828 11756
rect 17776 11713 17785 11747
rect 17785 11713 17819 11747
rect 17819 11713 17828 11747
rect 17776 11704 17828 11713
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 18972 11704 19024 11756
rect 22192 11704 22244 11756
rect 23664 11772 23716 11824
rect 25688 11772 25740 11824
rect 25964 11772 26016 11824
rect 23940 11704 23992 11756
rect 2596 11636 2648 11688
rect 4436 11636 4488 11688
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 5724 11636 5776 11688
rect 10140 11636 10192 11688
rect 14556 11636 14608 11688
rect 15752 11636 15804 11688
rect 17408 11636 17460 11688
rect 16120 11568 16172 11620
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 6644 11500 6696 11552
rect 7748 11500 7800 11552
rect 12440 11500 12492 11552
rect 13268 11500 13320 11552
rect 14648 11500 14700 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16856 11500 16908 11552
rect 17132 11500 17184 11552
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 17960 11568 18012 11620
rect 23848 11636 23900 11688
rect 27620 11704 27672 11756
rect 27896 11747 27948 11756
rect 27896 11713 27905 11747
rect 27905 11713 27939 11747
rect 27939 11713 27948 11747
rect 27896 11704 27948 11713
rect 27988 11747 28040 11756
rect 27988 11713 27997 11747
rect 27997 11713 28031 11747
rect 28031 11713 28040 11747
rect 27988 11704 28040 11713
rect 28080 11704 28132 11756
rect 29736 11772 29788 11824
rect 22560 11568 22612 11620
rect 27528 11636 27580 11688
rect 27804 11568 27856 11620
rect 28724 11568 28776 11620
rect 29644 11704 29696 11756
rect 29920 11636 29972 11688
rect 30196 11636 30248 11688
rect 29092 11568 29144 11620
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19064 11500 19116 11509
rect 22744 11500 22796 11552
rect 27344 11543 27396 11552
rect 27344 11509 27353 11543
rect 27353 11509 27387 11543
rect 27387 11509 27396 11543
rect 27344 11500 27396 11509
rect 31024 11500 31076 11552
rect 4871 11398 4923 11450
rect 4935 11398 4987 11450
rect 4999 11398 5051 11450
rect 5063 11398 5115 11450
rect 5127 11398 5179 11450
rect 12713 11398 12765 11450
rect 12777 11398 12829 11450
rect 12841 11398 12893 11450
rect 12905 11398 12957 11450
rect 12969 11398 13021 11450
rect 20555 11398 20607 11450
rect 20619 11398 20671 11450
rect 20683 11398 20735 11450
rect 20747 11398 20799 11450
rect 20811 11398 20863 11450
rect 28397 11398 28449 11450
rect 28461 11398 28513 11450
rect 28525 11398 28577 11450
rect 28589 11398 28641 11450
rect 28653 11398 28705 11450
rect 4712 11296 4764 11348
rect 6000 11296 6052 11348
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 6644 11228 6696 11280
rect 15292 11296 15344 11348
rect 17040 11296 17092 11348
rect 17408 11296 17460 11348
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 22376 11296 22428 11348
rect 23940 11296 23992 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 25872 11296 25924 11348
rect 13636 11228 13688 11280
rect 17776 11228 17828 11280
rect 5632 11160 5684 11212
rect 6000 11092 6052 11144
rect 2596 10956 2648 11008
rect 3424 10956 3476 11008
rect 5816 11024 5868 11076
rect 5908 11067 5960 11076
rect 5908 11033 5917 11067
rect 5917 11033 5951 11067
rect 5951 11033 5960 11067
rect 5908 11024 5960 11033
rect 6092 11024 6144 11076
rect 7564 11092 7616 11144
rect 8116 11092 8168 11144
rect 6828 11024 6880 11076
rect 7196 11024 7248 11076
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10232 11092 10284 11144
rect 15660 11160 15712 11212
rect 11060 11092 11112 11144
rect 11888 11092 11940 11144
rect 14372 11092 14424 11144
rect 14832 11092 14884 11144
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15568 11092 15620 11144
rect 18052 11160 18104 11212
rect 19064 11228 19116 11280
rect 17868 11092 17920 11144
rect 23756 11228 23808 11280
rect 20260 11092 20312 11144
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 23664 11160 23716 11212
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 10048 11024 10100 11076
rect 15476 11024 15528 11076
rect 15936 11024 15988 11076
rect 16948 11024 17000 11076
rect 8576 10999 8628 11008
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 14556 10956 14608 11008
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 17132 11024 17184 11076
rect 20168 11067 20220 11076
rect 20168 11033 20177 11067
rect 20177 11033 20211 11067
rect 20211 11033 20220 11067
rect 20168 11024 20220 11033
rect 23664 11024 23716 11076
rect 27436 11228 27488 11280
rect 30196 11339 30248 11348
rect 30196 11305 30205 11339
rect 30205 11305 30239 11339
rect 30239 11305 30248 11339
rect 30196 11296 30248 11305
rect 30748 11339 30800 11348
rect 30748 11305 30757 11339
rect 30757 11305 30791 11339
rect 30791 11305 30800 11339
rect 30748 11296 30800 11305
rect 30932 11339 30984 11348
rect 30932 11305 30941 11339
rect 30941 11305 30975 11339
rect 30975 11305 30984 11339
rect 30932 11296 30984 11305
rect 27620 11203 27672 11212
rect 27620 11169 27629 11203
rect 27629 11169 27663 11203
rect 27663 11169 27672 11203
rect 27620 11160 27672 11169
rect 29000 11160 29052 11212
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 25780 11092 25832 11101
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 27804 11092 27856 11144
rect 27988 11135 28040 11144
rect 27988 11101 27997 11135
rect 27997 11101 28031 11135
rect 28031 11101 28040 11135
rect 27988 11092 28040 11101
rect 17408 10956 17460 11008
rect 19616 10999 19668 11008
rect 19616 10965 19625 10999
rect 19625 10965 19659 10999
rect 19659 10965 19668 10999
rect 19616 10956 19668 10965
rect 24952 10956 25004 11008
rect 27528 11024 27580 11076
rect 28264 11024 28316 11076
rect 29184 11135 29236 11144
rect 29184 11101 29193 11135
rect 29193 11101 29227 11135
rect 29227 11101 29236 11135
rect 29184 11092 29236 11101
rect 29276 11024 29328 11076
rect 31944 11228 31996 11280
rect 31024 11203 31076 11212
rect 31024 11169 31033 11203
rect 31033 11169 31067 11203
rect 31067 11169 31076 11203
rect 31024 11160 31076 11169
rect 31300 11135 31352 11144
rect 31300 11101 31309 11135
rect 31309 11101 31343 11135
rect 31343 11101 31352 11135
rect 31300 11092 31352 11101
rect 30380 11024 30432 11076
rect 30748 11024 30800 11076
rect 26056 10999 26108 11008
rect 26056 10965 26065 10999
rect 26065 10965 26099 10999
rect 26099 10965 26108 10999
rect 26056 10956 26108 10965
rect 27620 10956 27672 11008
rect 27804 10999 27856 11008
rect 27804 10965 27813 10999
rect 27813 10965 27847 10999
rect 27847 10965 27856 10999
rect 27804 10956 27856 10965
rect 28724 10999 28776 11008
rect 28724 10965 28733 10999
rect 28733 10965 28767 10999
rect 28767 10965 28776 10999
rect 28724 10956 28776 10965
rect 8792 10854 8844 10906
rect 8856 10854 8908 10906
rect 8920 10854 8972 10906
rect 8984 10854 9036 10906
rect 9048 10854 9100 10906
rect 16634 10854 16686 10906
rect 16698 10854 16750 10906
rect 16762 10854 16814 10906
rect 16826 10854 16878 10906
rect 16890 10854 16942 10906
rect 24476 10854 24528 10906
rect 24540 10854 24592 10906
rect 24604 10854 24656 10906
rect 24668 10854 24720 10906
rect 24732 10854 24784 10906
rect 32318 10854 32370 10906
rect 32382 10854 32434 10906
rect 32446 10854 32498 10906
rect 32510 10854 32562 10906
rect 32574 10854 32626 10906
rect 3424 10752 3476 10804
rect 3976 10752 4028 10804
rect 10048 10795 10100 10804
rect 10048 10761 10057 10795
rect 10057 10761 10091 10795
rect 10091 10761 10100 10795
rect 10048 10752 10100 10761
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 13084 10684 13136 10736
rect 14464 10684 14516 10736
rect 14740 10727 14792 10736
rect 14740 10693 14749 10727
rect 14749 10693 14783 10727
rect 14783 10693 14792 10727
rect 14740 10684 14792 10693
rect 5724 10616 5776 10668
rect 6460 10616 6512 10668
rect 10232 10659 10284 10668
rect 10232 10625 10241 10659
rect 10241 10625 10275 10659
rect 10275 10625 10284 10659
rect 10232 10616 10284 10625
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 15292 10752 15344 10804
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 15384 10616 15436 10668
rect 15660 10752 15712 10804
rect 15844 10795 15896 10804
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 17960 10752 18012 10804
rect 18972 10752 19024 10804
rect 17224 10684 17276 10736
rect 2596 10591 2648 10600
rect 2596 10557 2605 10591
rect 2605 10557 2639 10591
rect 2639 10557 2648 10591
rect 2596 10548 2648 10557
rect 2688 10480 2740 10532
rect 9772 10548 9824 10600
rect 3424 10480 3476 10532
rect 8668 10480 8720 10532
rect 13728 10548 13780 10600
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 15752 10616 15804 10668
rect 13636 10480 13688 10532
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 17316 10548 17368 10600
rect 18236 10548 18288 10600
rect 18512 10616 18564 10668
rect 22008 10752 22060 10804
rect 23480 10752 23532 10804
rect 25596 10795 25648 10804
rect 25596 10761 25605 10795
rect 25605 10761 25639 10795
rect 25639 10761 25648 10795
rect 25596 10752 25648 10761
rect 27988 10752 28040 10804
rect 28816 10752 28868 10804
rect 19156 10727 19208 10736
rect 19156 10693 19165 10727
rect 19165 10693 19199 10727
rect 19199 10693 19208 10727
rect 19156 10684 19208 10693
rect 18788 10480 18840 10532
rect 5264 10412 5316 10464
rect 6828 10412 6880 10464
rect 9680 10412 9732 10464
rect 11796 10412 11848 10464
rect 13544 10412 13596 10464
rect 19800 10616 19852 10668
rect 19340 10548 19392 10600
rect 19524 10548 19576 10600
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 22560 10616 22612 10668
rect 23388 10727 23440 10736
rect 23388 10693 23397 10727
rect 23397 10693 23431 10727
rect 23431 10693 23440 10727
rect 23388 10684 23440 10693
rect 23296 10616 23348 10668
rect 26516 10684 26568 10736
rect 26608 10684 26660 10736
rect 29184 10684 29236 10736
rect 22468 10548 22520 10600
rect 21916 10480 21968 10532
rect 27344 10616 27396 10668
rect 27896 10616 27948 10668
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 28908 10659 28960 10668
rect 28908 10625 28917 10659
rect 28917 10625 28951 10659
rect 28951 10625 28960 10659
rect 28908 10616 28960 10625
rect 29736 10616 29788 10668
rect 31116 10752 31168 10804
rect 30104 10684 30156 10736
rect 30012 10659 30064 10668
rect 30012 10625 30021 10659
rect 30021 10625 30055 10659
rect 30055 10625 30064 10659
rect 30012 10616 30064 10625
rect 27988 10548 28040 10600
rect 28632 10548 28684 10600
rect 29000 10591 29052 10600
rect 29000 10557 29009 10591
rect 29009 10557 29043 10591
rect 29043 10557 29052 10591
rect 29000 10548 29052 10557
rect 30748 10659 30800 10668
rect 30748 10625 30757 10659
rect 30757 10625 30791 10659
rect 30791 10625 30800 10659
rect 30748 10616 30800 10625
rect 30564 10548 30616 10600
rect 31300 10616 31352 10668
rect 31760 10616 31812 10668
rect 26332 10480 26384 10532
rect 29276 10480 29328 10532
rect 20168 10412 20220 10464
rect 20352 10455 20404 10464
rect 20352 10421 20361 10455
rect 20361 10421 20395 10455
rect 20395 10421 20404 10455
rect 20352 10412 20404 10421
rect 22468 10412 22520 10464
rect 24400 10412 24452 10464
rect 27620 10412 27672 10464
rect 29644 10455 29696 10464
rect 29644 10421 29653 10455
rect 29653 10421 29687 10455
rect 29687 10421 29696 10455
rect 29644 10412 29696 10421
rect 29736 10412 29788 10464
rect 31024 10412 31076 10464
rect 4871 10310 4923 10362
rect 4935 10310 4987 10362
rect 4999 10310 5051 10362
rect 5063 10310 5115 10362
rect 5127 10310 5179 10362
rect 12713 10310 12765 10362
rect 12777 10310 12829 10362
rect 12841 10310 12893 10362
rect 12905 10310 12957 10362
rect 12969 10310 13021 10362
rect 20555 10310 20607 10362
rect 20619 10310 20671 10362
rect 20683 10310 20735 10362
rect 20747 10310 20799 10362
rect 20811 10310 20863 10362
rect 28397 10310 28449 10362
rect 28461 10310 28513 10362
rect 28525 10310 28577 10362
rect 28589 10310 28641 10362
rect 28653 10310 28705 10362
rect 2688 10251 2740 10260
rect 2688 10217 2697 10251
rect 2697 10217 2731 10251
rect 2731 10217 2740 10251
rect 2688 10208 2740 10217
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 3516 10208 3568 10260
rect 6092 10208 6144 10260
rect 10140 10208 10192 10260
rect 15292 10208 15344 10260
rect 15568 10208 15620 10260
rect 18420 10208 18472 10260
rect 18604 10208 18656 10260
rect 19524 10208 19576 10260
rect 19616 10208 19668 10260
rect 23112 10208 23164 10260
rect 23664 10208 23716 10260
rect 27620 10251 27672 10260
rect 27620 10217 27629 10251
rect 27629 10217 27663 10251
rect 27663 10217 27672 10251
rect 27620 10208 27672 10217
rect 31024 10251 31076 10260
rect 31024 10217 31033 10251
rect 31033 10217 31067 10251
rect 31067 10217 31076 10251
rect 31024 10208 31076 10217
rect 31760 10251 31812 10260
rect 31760 10217 31769 10251
rect 31769 10217 31803 10251
rect 31803 10217 31812 10251
rect 31760 10208 31812 10217
rect 3792 10140 3844 10192
rect 4160 10140 4212 10192
rect 15660 10140 15712 10192
rect 18512 10183 18564 10192
rect 18512 10149 18521 10183
rect 18521 10149 18555 10183
rect 18555 10149 18564 10183
rect 18512 10140 18564 10149
rect 18788 10140 18840 10192
rect 23204 10140 23256 10192
rect 3332 10004 3384 10056
rect 3608 10004 3660 10056
rect 3884 10004 3936 10056
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 6552 10047 6604 10056
rect 4620 10004 4672 10013
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 9680 10004 9732 10056
rect 11152 10004 11204 10056
rect 2872 9936 2924 9988
rect 5264 9936 5316 9988
rect 6828 9979 6880 9988
rect 6828 9945 6862 9979
rect 6862 9945 6880 9979
rect 6828 9936 6880 9945
rect 8576 9936 8628 9988
rect 11336 9979 11388 9988
rect 11336 9945 11370 9979
rect 11370 9945 11388 9979
rect 11336 9936 11388 9945
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 6736 9868 6788 9920
rect 11888 9868 11940 9920
rect 12532 9936 12584 9988
rect 13176 9979 13228 9988
rect 13176 9945 13185 9979
rect 13185 9945 13219 9979
rect 13219 9945 13228 9979
rect 13176 9936 13228 9945
rect 13728 9936 13780 9988
rect 15016 10072 15068 10124
rect 14924 10004 14976 10056
rect 17500 10072 17552 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 23388 10072 23440 10124
rect 15568 10047 15620 10056
rect 15108 9936 15160 9988
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 15016 9868 15068 9920
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 18328 10004 18380 10056
rect 20352 10004 20404 10056
rect 26792 10140 26844 10192
rect 27988 10140 28040 10192
rect 27804 10072 27856 10124
rect 29460 10072 29512 10124
rect 30012 10072 30064 10124
rect 30932 10115 30984 10124
rect 30932 10081 30941 10115
rect 30941 10081 30975 10115
rect 30975 10081 30984 10115
rect 30932 10072 30984 10081
rect 17316 9911 17368 9920
rect 17316 9877 17325 9911
rect 17325 9877 17359 9911
rect 17359 9877 17368 9911
rect 17316 9868 17368 9877
rect 17500 9911 17552 9920
rect 17500 9877 17527 9911
rect 17527 9877 17552 9911
rect 17500 9868 17552 9877
rect 18236 9936 18288 9988
rect 19248 9868 19300 9920
rect 23204 9979 23256 9988
rect 23204 9945 23213 9979
rect 23213 9945 23247 9979
rect 23247 9945 23256 9979
rect 23204 9936 23256 9945
rect 23664 9936 23716 9988
rect 24952 10047 25004 10056
rect 24952 10013 24994 10047
rect 24994 10013 25004 10047
rect 24952 10004 25004 10013
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 26056 10004 26108 10056
rect 26332 10047 26384 10056
rect 26332 10013 26341 10047
rect 26341 10013 26375 10047
rect 26375 10013 26384 10047
rect 26332 10004 26384 10013
rect 26516 10047 26568 10056
rect 26516 10013 26525 10047
rect 26525 10013 26559 10047
rect 26559 10013 26568 10047
rect 26516 10004 26568 10013
rect 26608 9936 26660 9988
rect 27436 10047 27488 10056
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 27712 10047 27764 10056
rect 27712 10013 27721 10047
rect 27721 10013 27755 10047
rect 27755 10013 27764 10047
rect 27712 10004 27764 10013
rect 28264 10004 28316 10056
rect 28724 10004 28776 10056
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 31116 10047 31168 10056
rect 31116 10013 31125 10047
rect 31125 10013 31159 10047
rect 31159 10013 31168 10047
rect 31116 10004 31168 10013
rect 19800 9911 19852 9920
rect 19800 9877 19809 9911
rect 19809 9877 19843 9911
rect 19843 9877 19852 9911
rect 19800 9868 19852 9877
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 25044 9911 25096 9920
rect 25044 9877 25053 9911
rect 25053 9877 25087 9911
rect 25087 9877 25096 9911
rect 25044 9868 25096 9877
rect 25964 9911 26016 9920
rect 25964 9877 25973 9911
rect 25973 9877 26007 9911
rect 26007 9877 26016 9911
rect 25964 9868 26016 9877
rect 27620 9868 27672 9920
rect 27988 9868 28040 9920
rect 30840 9979 30892 9988
rect 30840 9945 30849 9979
rect 30849 9945 30883 9979
rect 30883 9945 30892 9979
rect 30840 9936 30892 9945
rect 31944 10047 31996 10056
rect 31944 10013 31953 10047
rect 31953 10013 31987 10047
rect 31987 10013 31996 10047
rect 31944 10004 31996 10013
rect 8792 9766 8844 9818
rect 8856 9766 8908 9818
rect 8920 9766 8972 9818
rect 8984 9766 9036 9818
rect 9048 9766 9100 9818
rect 16634 9766 16686 9818
rect 16698 9766 16750 9818
rect 16762 9766 16814 9818
rect 16826 9766 16878 9818
rect 16890 9766 16942 9818
rect 24476 9766 24528 9818
rect 24540 9766 24592 9818
rect 24604 9766 24656 9818
rect 24668 9766 24720 9818
rect 24732 9766 24784 9818
rect 32318 9766 32370 9818
rect 32382 9766 32434 9818
rect 32446 9766 32498 9818
rect 32510 9766 32562 9818
rect 32574 9766 32626 9818
rect 2320 9664 2372 9716
rect 2228 9528 2280 9580
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 3056 9528 3108 9580
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 6092 9664 6144 9716
rect 6552 9664 6604 9716
rect 6368 9596 6420 9648
rect 14556 9664 14608 9716
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7012 9528 7064 9580
rect 12900 9596 12952 9648
rect 9680 9528 9732 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 11888 9571 11940 9580
rect 3056 9392 3108 9444
rect 5908 9460 5960 9512
rect 9956 9460 10008 9512
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 11336 9460 11388 9512
rect 12624 9528 12676 9580
rect 14464 9596 14516 9648
rect 15200 9639 15252 9648
rect 15200 9605 15209 9639
rect 15209 9605 15243 9639
rect 15243 9605 15252 9639
rect 15200 9596 15252 9605
rect 17132 9596 17184 9648
rect 17408 9596 17460 9648
rect 19340 9596 19392 9648
rect 19800 9664 19852 9716
rect 22192 9707 22244 9716
rect 22192 9673 22201 9707
rect 22201 9673 22235 9707
rect 22235 9673 22244 9707
rect 22192 9664 22244 9673
rect 25044 9664 25096 9716
rect 26056 9664 26108 9716
rect 19616 9596 19668 9648
rect 13084 9528 13136 9580
rect 13268 9571 13320 9580
rect 13268 9537 13302 9571
rect 13302 9537 13320 9571
rect 13268 9528 13320 9537
rect 12532 9460 12584 9512
rect 2964 9324 3016 9376
rect 3148 9324 3200 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 7564 9324 7616 9376
rect 15476 9528 15528 9580
rect 17316 9528 17368 9580
rect 18236 9528 18288 9580
rect 19248 9571 19300 9580
rect 19248 9537 19257 9571
rect 19257 9537 19291 9571
rect 19291 9537 19300 9571
rect 19248 9528 19300 9537
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 21916 9596 21968 9648
rect 22560 9596 22612 9648
rect 23664 9596 23716 9648
rect 25320 9639 25372 9648
rect 25320 9605 25329 9639
rect 25329 9605 25363 9639
rect 25363 9605 25372 9639
rect 25320 9596 25372 9605
rect 26148 9596 26200 9648
rect 26240 9639 26292 9648
rect 26240 9605 26249 9639
rect 26249 9605 26283 9639
rect 26283 9605 26292 9639
rect 26240 9596 26292 9605
rect 26608 9596 26660 9648
rect 26700 9596 26752 9648
rect 27252 9596 27304 9648
rect 15200 9460 15252 9512
rect 15384 9460 15436 9512
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 19340 9460 19392 9512
rect 20444 9460 20496 9512
rect 11612 9324 11664 9376
rect 11980 9324 12032 9376
rect 17316 9392 17368 9444
rect 18328 9392 18380 9444
rect 24308 9528 24360 9580
rect 27620 9571 27672 9580
rect 27620 9537 27629 9571
rect 27629 9537 27663 9571
rect 27663 9537 27672 9571
rect 27620 9528 27672 9537
rect 14740 9324 14792 9376
rect 17132 9324 17184 9376
rect 21088 9392 21140 9444
rect 21916 9392 21968 9444
rect 24952 9460 25004 9512
rect 27896 9707 27948 9716
rect 27896 9673 27905 9707
rect 27905 9673 27939 9707
rect 27939 9673 27948 9707
rect 27896 9664 27948 9673
rect 29460 9664 29512 9716
rect 30472 9664 30524 9716
rect 31116 9664 31168 9716
rect 28172 9528 28224 9580
rect 30840 9596 30892 9648
rect 19616 9324 19668 9376
rect 24768 9324 24820 9376
rect 26148 9392 26200 9444
rect 28816 9528 28868 9580
rect 29460 9571 29512 9580
rect 29460 9537 29469 9571
rect 29469 9537 29503 9571
rect 29503 9537 29512 9571
rect 29460 9528 29512 9537
rect 30288 9571 30340 9580
rect 30288 9537 30297 9571
rect 30297 9537 30331 9571
rect 30331 9537 30340 9571
rect 30288 9528 30340 9537
rect 29736 9460 29788 9512
rect 26240 9324 26292 9376
rect 26516 9324 26568 9376
rect 26792 9324 26844 9376
rect 27804 9324 27856 9376
rect 27896 9324 27948 9376
rect 29736 9324 29788 9376
rect 31484 9324 31536 9376
rect 4871 9222 4923 9274
rect 4935 9222 4987 9274
rect 4999 9222 5051 9274
rect 5063 9222 5115 9274
rect 5127 9222 5179 9274
rect 12713 9222 12765 9274
rect 12777 9222 12829 9274
rect 12841 9222 12893 9274
rect 12905 9222 12957 9274
rect 12969 9222 13021 9274
rect 20555 9222 20607 9274
rect 20619 9222 20671 9274
rect 20683 9222 20735 9274
rect 20747 9222 20799 9274
rect 20811 9222 20863 9274
rect 28397 9222 28449 9274
rect 28461 9222 28513 9274
rect 28525 9222 28577 9274
rect 28589 9222 28641 9274
rect 28653 9222 28705 9274
rect 4160 9120 4212 9172
rect 5724 9120 5776 9172
rect 6460 9120 6512 9172
rect 10232 9120 10284 9172
rect 12624 9120 12676 9172
rect 13176 9120 13228 9172
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 3240 9052 3292 9104
rect 3516 9052 3568 9104
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 2780 8916 2832 8968
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 3056 8984 3108 8993
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3700 8916 3752 8968
rect 7564 9052 7616 9104
rect 9128 9052 9180 9104
rect 9864 9052 9916 9104
rect 10876 9052 10928 9104
rect 13636 9052 13688 9104
rect 16028 9120 16080 9172
rect 7288 8984 7340 9036
rect 3332 8848 3384 8900
rect 4712 8916 4764 8968
rect 4620 8848 4672 8900
rect 5448 8891 5500 8900
rect 5448 8857 5457 8891
rect 5457 8857 5491 8891
rect 5491 8857 5500 8891
rect 5448 8848 5500 8857
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 6644 8848 6696 8900
rect 2964 8780 3016 8832
rect 3056 8780 3108 8832
rect 7656 8891 7708 8900
rect 7656 8857 7665 8891
rect 7665 8857 7699 8891
rect 7699 8857 7708 8891
rect 7656 8848 7708 8857
rect 8300 8916 8352 8968
rect 8484 8916 8536 8968
rect 9404 8916 9456 8968
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 11796 8959 11848 8968
rect 11796 8925 11814 8959
rect 11814 8925 11848 8959
rect 11796 8916 11848 8925
rect 11980 8916 12032 8968
rect 13084 8984 13136 9036
rect 12440 8916 12492 8968
rect 12716 8916 12768 8968
rect 13452 8916 13504 8968
rect 17592 9052 17644 9104
rect 18236 9120 18288 9172
rect 19340 9120 19392 9172
rect 19432 9120 19484 9172
rect 18512 9052 18564 9104
rect 14464 9027 14516 9036
rect 14464 8993 14473 9027
rect 14473 8993 14507 9027
rect 14507 8993 14516 9027
rect 14464 8984 14516 8993
rect 26608 9163 26660 9172
rect 26608 9129 26617 9163
rect 26617 9129 26651 9163
rect 26651 9129 26660 9163
rect 26608 9120 26660 9129
rect 26148 9052 26200 9104
rect 29000 9120 29052 9172
rect 14740 8959 14792 8968
rect 14740 8925 14774 8959
rect 14774 8925 14792 8959
rect 14740 8916 14792 8925
rect 15108 8916 15160 8968
rect 17040 8916 17092 8968
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 8116 8780 8168 8832
rect 12164 8848 12216 8900
rect 12348 8848 12400 8900
rect 10048 8780 10100 8832
rect 10232 8780 10284 8832
rect 17132 8848 17184 8900
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 20904 8916 20956 8968
rect 23480 8984 23532 9036
rect 19892 8848 19944 8900
rect 20444 8848 20496 8900
rect 21916 8916 21968 8968
rect 22468 8959 22520 8968
rect 22468 8925 22502 8959
rect 22502 8925 22520 8959
rect 22468 8916 22520 8925
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 21364 8848 21416 8900
rect 25964 8959 26016 8968
rect 25964 8925 25973 8959
rect 25973 8925 26007 8959
rect 26007 8925 26016 8959
rect 25964 8916 26016 8925
rect 26240 8916 26292 8968
rect 27712 8984 27764 9036
rect 28172 9027 28224 9036
rect 28172 8993 28181 9027
rect 28181 8993 28215 9027
rect 28215 8993 28224 9027
rect 28172 8984 28224 8993
rect 29644 8984 29696 9036
rect 26976 8916 27028 8968
rect 27804 8916 27856 8968
rect 28724 8916 28776 8968
rect 28908 8916 28960 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 16212 8780 16264 8832
rect 17224 8780 17276 8832
rect 18696 8823 18748 8832
rect 18696 8789 18721 8823
rect 18721 8789 18748 8823
rect 18696 8780 18748 8789
rect 19432 8780 19484 8832
rect 19616 8780 19668 8832
rect 22008 8780 22060 8832
rect 23664 8780 23716 8832
rect 25228 8780 25280 8832
rect 25780 8780 25832 8832
rect 27896 8780 27948 8832
rect 30380 8823 30432 8832
rect 30380 8789 30389 8823
rect 30389 8789 30423 8823
rect 30423 8789 30432 8823
rect 30380 8780 30432 8789
rect 8792 8678 8844 8730
rect 8856 8678 8908 8730
rect 8920 8678 8972 8730
rect 8984 8678 9036 8730
rect 9048 8678 9100 8730
rect 16634 8678 16686 8730
rect 16698 8678 16750 8730
rect 16762 8678 16814 8730
rect 16826 8678 16878 8730
rect 16890 8678 16942 8730
rect 24476 8678 24528 8730
rect 24540 8678 24592 8730
rect 24604 8678 24656 8730
rect 24668 8678 24720 8730
rect 24732 8678 24784 8730
rect 32318 8678 32370 8730
rect 32382 8678 32434 8730
rect 32446 8678 32498 8730
rect 32510 8678 32562 8730
rect 32574 8678 32626 8730
rect 3056 8576 3108 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 4620 8508 4672 8560
rect 8392 8576 8444 8628
rect 7288 8508 7340 8560
rect 8484 8508 8536 8560
rect 2044 8440 2096 8492
rect 2780 8440 2832 8492
rect 3332 8440 3384 8492
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 6000 8483 6052 8492
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 5540 8372 5592 8424
rect 2964 8304 3016 8356
rect 3792 8347 3844 8356
rect 3792 8313 3801 8347
rect 3801 8313 3835 8347
rect 3835 8313 3844 8347
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6368 8440 6420 8492
rect 7656 8440 7708 8492
rect 7932 8440 7984 8492
rect 10324 8576 10376 8628
rect 12532 8576 12584 8628
rect 13452 8576 13504 8628
rect 14648 8576 14700 8628
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 20260 8576 20312 8628
rect 22376 8619 22428 8628
rect 22376 8585 22385 8619
rect 22385 8585 22419 8619
rect 22419 8585 22428 8619
rect 22376 8576 22428 8585
rect 24308 8619 24360 8628
rect 24308 8585 24317 8619
rect 24317 8585 24351 8619
rect 24351 8585 24360 8619
rect 24308 8576 24360 8585
rect 24400 8576 24452 8628
rect 10232 8508 10284 8560
rect 10876 8508 10928 8560
rect 9956 8440 10008 8492
rect 11612 8508 11664 8560
rect 12348 8508 12400 8560
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 9772 8372 9824 8424
rect 12164 8440 12216 8492
rect 14464 8508 14516 8560
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 15108 8440 15160 8492
rect 16212 8440 16264 8492
rect 18512 8508 18564 8560
rect 21364 8508 21416 8560
rect 27620 8576 27672 8628
rect 29828 8576 29880 8628
rect 17500 8483 17552 8492
rect 17500 8449 17534 8483
rect 17534 8449 17552 8483
rect 17500 8440 17552 8449
rect 18696 8440 18748 8492
rect 20720 8440 20772 8492
rect 21180 8440 21232 8492
rect 21916 8440 21968 8492
rect 23480 8483 23532 8492
rect 23480 8449 23498 8483
rect 23498 8449 23532 8483
rect 23480 8440 23532 8449
rect 12624 8372 12676 8424
rect 3792 8304 3844 8313
rect 5724 8236 5776 8288
rect 6644 8236 6696 8288
rect 7104 8304 7156 8356
rect 11612 8304 11664 8356
rect 11704 8347 11756 8356
rect 11704 8313 11713 8347
rect 11713 8313 11747 8347
rect 11747 8313 11756 8347
rect 11704 8304 11756 8313
rect 14556 8304 14608 8356
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 10324 8236 10376 8245
rect 10968 8236 11020 8288
rect 14648 8236 14700 8288
rect 17224 8236 17276 8288
rect 23572 8236 23624 8288
rect 24860 8440 24912 8492
rect 25412 8483 25464 8492
rect 25412 8449 25446 8483
rect 25446 8449 25464 8483
rect 25412 8440 25464 8449
rect 27252 8440 27304 8492
rect 30288 8508 30340 8560
rect 30380 8440 30432 8492
rect 24768 8236 24820 8288
rect 27804 8236 27856 8288
rect 4871 8134 4923 8186
rect 4935 8134 4987 8186
rect 4999 8134 5051 8186
rect 5063 8134 5115 8186
rect 5127 8134 5179 8186
rect 12713 8134 12765 8186
rect 12777 8134 12829 8186
rect 12841 8134 12893 8186
rect 12905 8134 12957 8186
rect 12969 8134 13021 8186
rect 20555 8134 20607 8186
rect 20619 8134 20671 8186
rect 20683 8134 20735 8186
rect 20747 8134 20799 8186
rect 20811 8134 20863 8186
rect 28397 8134 28449 8186
rect 28461 8134 28513 8186
rect 28525 8134 28577 8186
rect 28589 8134 28641 8186
rect 28653 8134 28705 8186
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 7012 8032 7064 8084
rect 8300 8032 8352 8084
rect 9496 8032 9548 8084
rect 17040 8032 17092 8084
rect 17500 8032 17552 8084
rect 19892 8075 19944 8084
rect 19892 8041 19901 8075
rect 19901 8041 19935 8075
rect 19935 8041 19944 8075
rect 19892 8032 19944 8041
rect 10232 8007 10284 8016
rect 10232 7973 10241 8007
rect 10241 7973 10275 8007
rect 10275 7973 10284 8007
rect 10232 7964 10284 7973
rect 17408 7964 17460 8016
rect 6920 7896 6972 7948
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 17040 7896 17092 7948
rect 2872 7828 2924 7880
rect 3240 7828 3292 7880
rect 7104 7828 7156 7880
rect 9956 7871 10008 7880
rect 6368 7760 6420 7812
rect 7012 7760 7064 7812
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 11060 7828 11112 7880
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 11888 7828 11940 7880
rect 14556 7828 14608 7880
rect 17132 7828 17184 7880
rect 17316 7828 17368 7880
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 17868 7828 17920 7880
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 19616 7828 19668 7880
rect 21180 8075 21232 8084
rect 21180 8041 21189 8075
rect 21189 8041 21223 8075
rect 21223 8041 21232 8075
rect 21180 8032 21232 8041
rect 23572 8032 23624 8084
rect 24308 8032 24360 8084
rect 25412 8075 25464 8084
rect 25412 8041 25421 8075
rect 25421 8041 25455 8075
rect 25455 8041 25464 8075
rect 25412 8032 25464 8041
rect 27252 8032 27304 8084
rect 28172 8032 28224 8084
rect 22376 7896 22428 7948
rect 22560 7896 22612 7948
rect 23480 7964 23532 8016
rect 27804 7896 27856 7948
rect 2872 7692 2924 7744
rect 3884 7692 3936 7744
rect 5264 7692 5316 7744
rect 6736 7692 6788 7744
rect 7196 7692 7248 7744
rect 8668 7692 8720 7744
rect 9404 7692 9456 7744
rect 10140 7760 10192 7812
rect 15384 7760 15436 7812
rect 16396 7803 16448 7812
rect 16396 7769 16405 7803
rect 16405 7769 16439 7803
rect 16439 7769 16448 7803
rect 16396 7760 16448 7769
rect 17684 7760 17736 7812
rect 9588 7692 9640 7744
rect 13176 7735 13228 7744
rect 13176 7701 13185 7735
rect 13185 7701 13219 7735
rect 13219 7701 13228 7735
rect 13176 7692 13228 7701
rect 13728 7692 13780 7744
rect 13820 7692 13872 7744
rect 15936 7692 15988 7744
rect 20260 7692 20312 7744
rect 22376 7760 22428 7812
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 25228 7871 25280 7880
rect 25228 7837 25237 7871
rect 25237 7837 25271 7871
rect 25271 7837 25280 7871
rect 25228 7828 25280 7837
rect 26792 7871 26844 7880
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 27620 7871 27672 7880
rect 27620 7837 27629 7871
rect 27629 7837 27663 7871
rect 27663 7837 27672 7871
rect 27620 7828 27672 7837
rect 23296 7760 23348 7812
rect 24400 7692 24452 7744
rect 8792 7590 8844 7642
rect 8856 7590 8908 7642
rect 8920 7590 8972 7642
rect 8984 7590 9036 7642
rect 9048 7590 9100 7642
rect 16634 7590 16686 7642
rect 16698 7590 16750 7642
rect 16762 7590 16814 7642
rect 16826 7590 16878 7642
rect 16890 7590 16942 7642
rect 24476 7590 24528 7642
rect 24540 7590 24592 7642
rect 24604 7590 24656 7642
rect 24668 7590 24720 7642
rect 24732 7590 24784 7642
rect 32318 7590 32370 7642
rect 32382 7590 32434 7642
rect 32446 7590 32498 7642
rect 32510 7590 32562 7642
rect 32574 7590 32626 7642
rect 2964 7488 3016 7540
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 2872 7352 2924 7404
rect 5632 7488 5684 7540
rect 7012 7488 7064 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 9496 7531 9548 7540
rect 9496 7497 9505 7531
rect 9505 7497 9539 7531
rect 9539 7497 9548 7531
rect 9496 7488 9548 7497
rect 6644 7420 6696 7472
rect 5724 7352 5776 7404
rect 3240 7284 3292 7336
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 5540 7284 5592 7336
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 8668 7420 8720 7472
rect 9404 7420 9456 7472
rect 9588 7420 9640 7472
rect 10140 7463 10192 7472
rect 10140 7429 10165 7463
rect 10165 7429 10192 7463
rect 10140 7420 10192 7429
rect 8300 7352 8352 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 9772 7352 9824 7404
rect 10324 7352 10376 7404
rect 11336 7488 11388 7540
rect 12256 7488 12308 7540
rect 10968 7420 11020 7472
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 16396 7488 16448 7540
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 19524 7488 19576 7540
rect 21640 7488 21692 7540
rect 12256 7395 12308 7404
rect 3332 7216 3384 7268
rect 4252 7216 4304 7268
rect 9588 7284 9640 7336
rect 12256 7361 12298 7395
rect 12298 7361 12308 7395
rect 12256 7352 12308 7361
rect 13176 7352 13228 7404
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 11612 7284 11664 7336
rect 8116 7216 8168 7268
rect 9956 7216 10008 7268
rect 4436 7148 4488 7200
rect 6552 7148 6604 7200
rect 8576 7191 8628 7200
rect 8576 7157 8585 7191
rect 8585 7157 8619 7191
rect 8619 7157 8628 7191
rect 8576 7148 8628 7157
rect 13084 7284 13136 7336
rect 13452 7216 13504 7268
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 18604 7352 18656 7404
rect 22652 7420 22704 7472
rect 24308 7531 24360 7540
rect 24308 7497 24317 7531
rect 24317 7497 24351 7531
rect 24351 7497 24360 7531
rect 24308 7488 24360 7497
rect 24400 7488 24452 7540
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 20444 7284 20496 7336
rect 23020 7284 23072 7336
rect 24584 7352 24636 7404
rect 24860 7352 24912 7404
rect 10416 7148 10468 7200
rect 17960 7216 18012 7268
rect 20260 7216 20312 7268
rect 22468 7216 22520 7268
rect 17132 7148 17184 7200
rect 20444 7148 20496 7200
rect 21180 7148 21232 7200
rect 21732 7148 21784 7200
rect 23664 7216 23716 7268
rect 24584 7216 24636 7268
rect 24676 7216 24728 7268
rect 4871 7046 4923 7098
rect 4935 7046 4987 7098
rect 4999 7046 5051 7098
rect 5063 7046 5115 7098
rect 5127 7046 5179 7098
rect 12713 7046 12765 7098
rect 12777 7046 12829 7098
rect 12841 7046 12893 7098
rect 12905 7046 12957 7098
rect 12969 7046 13021 7098
rect 20555 7046 20607 7098
rect 20619 7046 20671 7098
rect 20683 7046 20735 7098
rect 20747 7046 20799 7098
rect 20811 7046 20863 7098
rect 28397 7046 28449 7098
rect 28461 7046 28513 7098
rect 28525 7046 28577 7098
rect 28589 7046 28641 7098
rect 28653 7046 28705 7098
rect 4252 6944 4304 6996
rect 5356 6944 5408 6996
rect 5540 6944 5592 6996
rect 6368 6944 6420 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 3056 6919 3108 6928
rect 3056 6885 3065 6919
rect 3065 6885 3099 6919
rect 3099 6885 3108 6919
rect 3056 6876 3108 6885
rect 3792 6808 3844 6860
rect 2688 6740 2740 6792
rect 3332 6740 3384 6792
rect 3976 6740 4028 6792
rect 4344 6740 4396 6792
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5264 6740 5316 6792
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7748 6740 7800 6792
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8576 6808 8628 6860
rect 9404 6851 9456 6860
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 9680 6808 9732 6860
rect 9496 6740 9548 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 12256 6851 12308 6860
rect 12256 6817 12265 6851
rect 12265 6817 12299 6851
rect 12299 6817 12308 6851
rect 12256 6808 12308 6817
rect 12440 6808 12492 6860
rect 13820 6876 13872 6928
rect 14832 6808 14884 6860
rect 17224 6944 17276 6996
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 20444 6987 20496 6996
rect 20444 6953 20453 6987
rect 20453 6953 20487 6987
rect 20487 6953 20496 6987
rect 20444 6944 20496 6953
rect 20812 6876 20864 6928
rect 21364 6876 21416 6928
rect 21732 6876 21784 6928
rect 16120 6808 16172 6860
rect 17316 6808 17368 6860
rect 17592 6808 17644 6860
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 12164 6783 12216 6792
rect 12164 6749 12173 6783
rect 12173 6749 12207 6783
rect 12207 6749 12216 6783
rect 12164 6740 12216 6749
rect 15844 6740 15896 6792
rect 16948 6740 17000 6792
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 17224 6740 17276 6792
rect 19616 6740 19668 6792
rect 20352 6740 20404 6792
rect 24676 6944 24728 6996
rect 22376 6919 22428 6928
rect 22376 6885 22385 6919
rect 22385 6885 22419 6919
rect 22419 6885 22428 6919
rect 22376 6876 22428 6885
rect 22560 6808 22612 6860
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 21088 6740 21140 6792
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 21732 6783 21784 6792
rect 21732 6749 21741 6783
rect 21741 6749 21775 6783
rect 21775 6749 21784 6783
rect 21732 6740 21784 6749
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 9772 6604 9824 6656
rect 11980 6604 12032 6656
rect 12440 6604 12492 6656
rect 18144 6604 18196 6656
rect 20076 6604 20128 6656
rect 21088 6604 21140 6656
rect 21824 6604 21876 6656
rect 23020 6740 23072 6792
rect 23296 6604 23348 6656
rect 8792 6502 8844 6554
rect 8856 6502 8908 6554
rect 8920 6502 8972 6554
rect 8984 6502 9036 6554
rect 9048 6502 9100 6554
rect 16634 6502 16686 6554
rect 16698 6502 16750 6554
rect 16762 6502 16814 6554
rect 16826 6502 16878 6554
rect 16890 6502 16942 6554
rect 24476 6502 24528 6554
rect 24540 6502 24592 6554
rect 24604 6502 24656 6554
rect 24668 6502 24720 6554
rect 24732 6502 24784 6554
rect 32318 6502 32370 6554
rect 32382 6502 32434 6554
rect 32446 6502 32498 6554
rect 32510 6502 32562 6554
rect 32574 6502 32626 6554
rect 4160 6400 4212 6452
rect 4620 6400 4672 6452
rect 4344 6375 4396 6384
rect 4344 6341 4353 6375
rect 4353 6341 4387 6375
rect 4387 6341 4396 6375
rect 10140 6400 10192 6452
rect 13728 6400 13780 6452
rect 17132 6400 17184 6452
rect 20076 6443 20128 6452
rect 20076 6409 20085 6443
rect 20085 6409 20119 6443
rect 20119 6409 20128 6443
rect 20076 6400 20128 6409
rect 21548 6400 21600 6452
rect 4344 6332 4396 6341
rect 5264 6375 5316 6384
rect 5264 6341 5273 6375
rect 5273 6341 5307 6375
rect 5307 6341 5316 6375
rect 5264 6332 5316 6341
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 4988 6264 5040 6316
rect 8300 6264 8352 6316
rect 8116 6196 8168 6248
rect 8576 6264 8628 6316
rect 11520 6332 11572 6384
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 14832 6264 14884 6316
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 16488 6264 16540 6316
rect 17316 6264 17368 6316
rect 19616 6375 19668 6384
rect 19616 6341 19625 6375
rect 19625 6341 19659 6375
rect 19659 6341 19668 6375
rect 19616 6332 19668 6341
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 12440 6060 12492 6112
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 17500 6239 17552 6248
rect 17500 6205 17509 6239
rect 17509 6205 17543 6239
rect 17543 6205 17552 6239
rect 17500 6196 17552 6205
rect 17224 6128 17276 6180
rect 16212 6060 16264 6112
rect 16488 6060 16540 6112
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 18604 6264 18656 6316
rect 19340 6128 19392 6180
rect 20260 6128 20312 6180
rect 20444 6128 20496 6180
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 21088 6307 21140 6316
rect 21088 6273 21104 6307
rect 21104 6273 21140 6307
rect 21088 6264 21140 6273
rect 21180 6307 21232 6316
rect 21180 6273 21189 6307
rect 21189 6273 21223 6307
rect 21223 6273 21232 6307
rect 21180 6264 21232 6273
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 21456 6196 21508 6248
rect 21732 6196 21784 6248
rect 20904 6128 20956 6180
rect 4871 5958 4923 6010
rect 4935 5958 4987 6010
rect 4999 5958 5051 6010
rect 5063 5958 5115 6010
rect 5127 5958 5179 6010
rect 12713 5958 12765 6010
rect 12777 5958 12829 6010
rect 12841 5958 12893 6010
rect 12905 5958 12957 6010
rect 12969 5958 13021 6010
rect 20555 5958 20607 6010
rect 20619 5958 20671 6010
rect 20683 5958 20735 6010
rect 20747 5958 20799 6010
rect 20811 5958 20863 6010
rect 28397 5958 28449 6010
rect 28461 5958 28513 6010
rect 28525 5958 28577 6010
rect 28589 5958 28641 6010
rect 28653 5958 28705 6010
rect 11980 5856 12032 5908
rect 13176 5856 13228 5908
rect 17132 5899 17184 5908
rect 17132 5865 17141 5899
rect 17141 5865 17175 5899
rect 17175 5865 17184 5899
rect 17132 5856 17184 5865
rect 18604 5856 18656 5908
rect 20996 5856 21048 5908
rect 21088 5856 21140 5908
rect 21640 5899 21692 5908
rect 21640 5865 21649 5899
rect 21649 5865 21683 5899
rect 21683 5865 21692 5899
rect 21640 5856 21692 5865
rect 22468 5899 22520 5908
rect 22468 5865 22477 5899
rect 22477 5865 22511 5899
rect 22511 5865 22520 5899
rect 22468 5856 22520 5865
rect 13820 5788 13872 5840
rect 18144 5788 18196 5840
rect 20444 5788 20496 5840
rect 16212 5763 16264 5772
rect 16212 5729 16221 5763
rect 16221 5729 16255 5763
rect 16255 5729 16264 5763
rect 16212 5720 16264 5729
rect 17500 5720 17552 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 12164 5652 12216 5704
rect 14832 5652 14884 5704
rect 17224 5652 17276 5704
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 21088 5720 21140 5772
rect 21548 5788 21600 5840
rect 21824 5652 21876 5704
rect 23020 5652 23072 5704
rect 17132 5584 17184 5636
rect 17316 5516 17368 5568
rect 21732 5516 21784 5568
rect 8792 5414 8844 5466
rect 8856 5414 8908 5466
rect 8920 5414 8972 5466
rect 8984 5414 9036 5466
rect 9048 5414 9100 5466
rect 16634 5414 16686 5466
rect 16698 5414 16750 5466
rect 16762 5414 16814 5466
rect 16826 5414 16878 5466
rect 16890 5414 16942 5466
rect 24476 5414 24528 5466
rect 24540 5414 24592 5466
rect 24604 5414 24656 5466
rect 24668 5414 24720 5466
rect 24732 5414 24784 5466
rect 32318 5414 32370 5466
rect 32382 5414 32434 5466
rect 32446 5414 32498 5466
rect 32510 5414 32562 5466
rect 32574 5414 32626 5466
rect 17040 5355 17092 5364
rect 17040 5321 17049 5355
rect 17049 5321 17083 5355
rect 17083 5321 17092 5355
rect 17040 5312 17092 5321
rect 20904 5312 20956 5364
rect 21824 5312 21876 5364
rect 17132 5244 17184 5296
rect 21732 5244 21784 5296
rect 17500 5176 17552 5228
rect 19616 5176 19668 5228
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 21364 5219 21416 5228
rect 21364 5185 21373 5219
rect 21373 5185 21407 5219
rect 21407 5185 21416 5219
rect 21364 5176 21416 5185
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 4871 4870 4923 4922
rect 4935 4870 4987 4922
rect 4999 4870 5051 4922
rect 5063 4870 5115 4922
rect 5127 4870 5179 4922
rect 12713 4870 12765 4922
rect 12777 4870 12829 4922
rect 12841 4870 12893 4922
rect 12905 4870 12957 4922
rect 12969 4870 13021 4922
rect 20555 4870 20607 4922
rect 20619 4870 20671 4922
rect 20683 4870 20735 4922
rect 20747 4870 20799 4922
rect 20811 4870 20863 4922
rect 28397 4870 28449 4922
rect 28461 4870 28513 4922
rect 28525 4870 28577 4922
rect 28589 4870 28641 4922
rect 28653 4870 28705 4922
rect 8792 4326 8844 4378
rect 8856 4326 8908 4378
rect 8920 4326 8972 4378
rect 8984 4326 9036 4378
rect 9048 4326 9100 4378
rect 16634 4326 16686 4378
rect 16698 4326 16750 4378
rect 16762 4326 16814 4378
rect 16826 4326 16878 4378
rect 16890 4326 16942 4378
rect 24476 4326 24528 4378
rect 24540 4326 24592 4378
rect 24604 4326 24656 4378
rect 24668 4326 24720 4378
rect 24732 4326 24784 4378
rect 32318 4326 32370 4378
rect 32382 4326 32434 4378
rect 32446 4326 32498 4378
rect 32510 4326 32562 4378
rect 32574 4326 32626 4378
rect 4871 3782 4923 3834
rect 4935 3782 4987 3834
rect 4999 3782 5051 3834
rect 5063 3782 5115 3834
rect 5127 3782 5179 3834
rect 12713 3782 12765 3834
rect 12777 3782 12829 3834
rect 12841 3782 12893 3834
rect 12905 3782 12957 3834
rect 12969 3782 13021 3834
rect 20555 3782 20607 3834
rect 20619 3782 20671 3834
rect 20683 3782 20735 3834
rect 20747 3782 20799 3834
rect 20811 3782 20863 3834
rect 28397 3782 28449 3834
rect 28461 3782 28513 3834
rect 28525 3782 28577 3834
rect 28589 3782 28641 3834
rect 28653 3782 28705 3834
rect 8792 3238 8844 3290
rect 8856 3238 8908 3290
rect 8920 3238 8972 3290
rect 8984 3238 9036 3290
rect 9048 3238 9100 3290
rect 16634 3238 16686 3290
rect 16698 3238 16750 3290
rect 16762 3238 16814 3290
rect 16826 3238 16878 3290
rect 16890 3238 16942 3290
rect 24476 3238 24528 3290
rect 24540 3238 24592 3290
rect 24604 3238 24656 3290
rect 24668 3238 24720 3290
rect 24732 3238 24784 3290
rect 32318 3238 32370 3290
rect 32382 3238 32434 3290
rect 32446 3238 32498 3290
rect 32510 3238 32562 3290
rect 32574 3238 32626 3290
rect 4871 2694 4923 2746
rect 4935 2694 4987 2746
rect 4999 2694 5051 2746
rect 5063 2694 5115 2746
rect 5127 2694 5179 2746
rect 12713 2694 12765 2746
rect 12777 2694 12829 2746
rect 12841 2694 12893 2746
rect 12905 2694 12957 2746
rect 12969 2694 13021 2746
rect 20555 2694 20607 2746
rect 20619 2694 20671 2746
rect 20683 2694 20735 2746
rect 20747 2694 20799 2746
rect 20811 2694 20863 2746
rect 28397 2694 28449 2746
rect 28461 2694 28513 2746
rect 28525 2694 28577 2746
rect 28589 2694 28641 2746
rect 28653 2694 28705 2746
rect 8792 2150 8844 2202
rect 8856 2150 8908 2202
rect 8920 2150 8972 2202
rect 8984 2150 9036 2202
rect 9048 2150 9100 2202
rect 16634 2150 16686 2202
rect 16698 2150 16750 2202
rect 16762 2150 16814 2202
rect 16826 2150 16878 2202
rect 16890 2150 16942 2202
rect 24476 2150 24528 2202
rect 24540 2150 24592 2202
rect 24604 2150 24656 2202
rect 24668 2150 24720 2202
rect 24732 2150 24784 2202
rect 32318 2150 32370 2202
rect 32382 2150 32434 2202
rect 32446 2150 32498 2202
rect 32510 2150 32562 2202
rect 32574 2150 32626 2202
rect 4871 1606 4923 1658
rect 4935 1606 4987 1658
rect 4999 1606 5051 1658
rect 5063 1606 5115 1658
rect 5127 1606 5179 1658
rect 12713 1606 12765 1658
rect 12777 1606 12829 1658
rect 12841 1606 12893 1658
rect 12905 1606 12957 1658
rect 12969 1606 13021 1658
rect 20555 1606 20607 1658
rect 20619 1606 20671 1658
rect 20683 1606 20735 1658
rect 20747 1606 20799 1658
rect 20811 1606 20863 1658
rect 28397 1606 28449 1658
rect 28461 1606 28513 1658
rect 28525 1606 28577 1658
rect 28589 1606 28641 1658
rect 28653 1606 28705 1658
rect 8792 1062 8844 1114
rect 8856 1062 8908 1114
rect 8920 1062 8972 1114
rect 8984 1062 9036 1114
rect 9048 1062 9100 1114
rect 16634 1062 16686 1114
rect 16698 1062 16750 1114
rect 16762 1062 16814 1114
rect 16826 1062 16878 1114
rect 16890 1062 16942 1114
rect 24476 1062 24528 1114
rect 24540 1062 24592 1114
rect 24604 1062 24656 1114
rect 24668 1062 24720 1114
rect 24732 1062 24784 1114
rect 32318 1062 32370 1114
rect 32382 1062 32434 1114
rect 32446 1062 32498 1114
rect 32510 1062 32562 1114
rect 32574 1062 32626 1114
<< metal2 >>
rect 2962 21448 3018 21457
rect 2962 21383 3018 21392
rect 4434 21448 4490 21457
rect 4434 21383 4490 21392
rect 4802 21448 4858 21457
rect 4802 21383 4858 21392
rect 5538 21448 5594 21457
rect 5538 21383 5594 21392
rect 6090 21448 6146 21457
rect 6090 21383 6146 21392
rect 8206 21448 8262 21457
rect 8206 21383 8262 21392
rect 9678 21448 9734 21457
rect 9678 21383 9734 21392
rect 11794 21448 11850 21457
rect 11794 21383 11850 21392
rect 13818 21448 13874 21457
rect 13818 21383 13874 21392
rect 14186 21448 14242 21457
rect 14186 21383 14242 21392
rect 15842 21448 15898 21457
rect 15842 21383 15898 21392
rect 28262 21448 28318 21457
rect 28262 21383 28318 21392
rect 28722 21448 28778 21457
rect 28722 21383 28778 21392
rect 29458 21448 29514 21457
rect 29458 21383 29514 21392
rect 31666 21448 31722 21457
rect 31722 21406 31892 21434
rect 31666 21383 31722 21392
rect 2976 19922 3004 21383
rect 4448 20602 4476 21383
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4816 20534 4844 21383
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4908 20602 4936 20742
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4724 20058 4752 20402
rect 4871 20156 5179 20165
rect 4871 20154 4877 20156
rect 4933 20154 4957 20156
rect 5013 20154 5037 20156
rect 5093 20154 5117 20156
rect 5173 20154 5179 20156
rect 4933 20102 4935 20154
rect 5115 20102 5117 20154
rect 4871 20100 4877 20102
rect 4933 20100 4957 20102
rect 5013 20100 5037 20102
rect 5093 20100 5117 20102
rect 5173 20100 5179 20102
rect 4871 20091 5179 20100
rect 5368 20058 5396 20810
rect 5552 20398 5580 21383
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 4068 19848 4120 19854
rect 4120 19808 4200 19836
rect 4068 19790 4120 19796
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 1766 19544 1822 19553
rect 1766 19479 1768 19488
rect 1820 19479 1822 19488
rect 1768 19450 1820 19456
rect 2792 19446 2820 19654
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 2240 18902 2268 19314
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18086 2176 18702
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2240 18086 2268 18566
rect 2608 18426 2636 18906
rect 2884 18630 2912 19246
rect 2976 18766 3004 19246
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1596 16250 1624 17847
rect 2148 17610 2176 18022
rect 2424 17882 2452 18294
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2056 16998 2084 17478
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16590 2084 16934
rect 2148 16590 2176 17546
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 2056 16114 2084 16526
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 16182 2360 16458
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2148 13326 2176 15302
rect 2424 14414 2452 17818
rect 2700 17202 2728 18158
rect 3068 17882 3096 18226
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3160 17746 3188 19314
rect 3252 18426 3280 19790
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3528 19514 3556 19722
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3436 18766 3464 19314
rect 4172 19310 4200 19808
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3068 17270 3096 17614
rect 3148 17604 3200 17610
rect 3200 17564 3280 17592
rect 3148 17546 3200 17552
rect 3056 17264 3108 17270
rect 3108 17212 3188 17218
rect 3056 17206 3188 17212
rect 2688 17196 2740 17202
rect 3068 17190 3188 17206
rect 3252 17202 3280 17564
rect 3344 17338 3372 18158
rect 3436 17814 3464 18702
rect 3514 17912 3570 17921
rect 3988 17882 4016 19246
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 4080 18630 4108 18838
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 3514 17847 3570 17856
rect 3608 17876 3660 17882
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 2688 17138 2740 17144
rect 2700 16658 2728 17138
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3068 16658 3096 16934
rect 3160 16658 3188 17190
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3252 16658 3280 17138
rect 3344 17066 3372 17274
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3436 16998 3464 17274
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2884 16250 2912 16390
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2240 12850 2268 13670
rect 2424 13258 2452 13670
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2424 12850 2452 13194
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2608 11694 2636 14894
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2700 12986 2728 13262
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2884 12850 2912 15574
rect 3068 15026 3096 16594
rect 3252 15502 3280 16594
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3528 15434 3556 17847
rect 3608 17818 3660 17824
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3620 17338 3648 17818
rect 3988 17678 4016 17818
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3620 15978 3648 16526
rect 3804 16114 3832 17478
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15638 3648 15914
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3804 15502 3832 16050
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 13530 3096 14214
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3068 13326 3096 13466
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12714 2912 12786
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2976 11898 3004 13262
rect 3160 13138 3188 14554
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 13938 3464 14214
rect 3528 14074 3556 14282
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3528 13938 3556 14010
rect 3620 13938 3648 15302
rect 3988 15026 4016 17614
rect 4080 16182 4108 18566
rect 4172 18222 4200 19246
rect 4356 18970 4384 19654
rect 4871 19068 5179 19077
rect 4871 19066 4877 19068
rect 4933 19066 4957 19068
rect 5013 19066 5037 19068
rect 5093 19066 5117 19068
rect 5173 19066 5179 19068
rect 4933 19014 4935 19066
rect 5115 19014 5117 19066
rect 4871 19012 4877 19014
rect 4933 19012 4957 19014
rect 5013 19012 5037 19014
rect 5093 19012 5117 19014
rect 5173 19012 5179 19014
rect 4871 19003 5179 19012
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 5368 18358 5396 19994
rect 5828 19242 5856 20402
rect 6012 20058 6040 20402
rect 6104 20330 6132 21383
rect 8114 20632 8170 20641
rect 8114 20567 8116 20576
rect 8168 20567 8170 20576
rect 8116 20538 8168 20544
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6564 19514 6592 20402
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6840 19378 6868 20198
rect 8128 19938 8156 20198
rect 8220 20058 8248 21383
rect 9494 20904 9550 20913
rect 9494 20839 9550 20848
rect 8792 20700 9100 20709
rect 8792 20698 8798 20700
rect 8854 20698 8878 20700
rect 8934 20698 8958 20700
rect 9014 20698 9038 20700
rect 9094 20698 9100 20700
rect 8854 20646 8856 20698
rect 9036 20646 9038 20698
rect 8792 20644 8798 20646
rect 8854 20644 8878 20646
rect 8934 20644 8958 20646
rect 9014 20644 9038 20646
rect 9094 20644 9100 20646
rect 8792 20635 9100 20644
rect 9508 20602 9536 20839
rect 9692 20602 9720 21383
rect 11058 21312 11114 21321
rect 11058 21247 11114 21256
rect 11702 21312 11758 21321
rect 11702 21247 11758 21256
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8576 19984 8628 19990
rect 8128 19922 8248 19938
rect 8576 19926 8628 19932
rect 8128 19916 8260 19922
rect 8128 19910 8208 19916
rect 8208 19858 8260 19864
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5828 18834 5856 19178
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 6932 18426 6960 19110
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4172 17202 4200 18158
rect 4448 17882 4476 18226
rect 7024 18154 7052 19790
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7116 18970 7144 19314
rect 8036 19242 8064 19314
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18222 7144 18566
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7208 18086 7236 19110
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 4871 17980 5179 17989
rect 4871 17978 4877 17980
rect 4933 17978 4957 17980
rect 5013 17978 5037 17980
rect 5093 17978 5117 17980
rect 5173 17978 5179 17980
rect 4933 17926 4935 17978
rect 5115 17926 5117 17978
rect 4871 17924 4877 17926
rect 4933 17924 4957 17926
rect 5013 17924 5037 17926
rect 5093 17924 5117 17926
rect 5173 17924 5179 17926
rect 4871 17915 5179 17924
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4172 16794 4200 17138
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4264 16250 4292 16458
rect 4356 16454 4384 17138
rect 5368 17066 5396 17478
rect 5552 17338 5580 17614
rect 6104 17610 6132 18022
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 6104 17202 6132 17546
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6012 17082 6040 17138
rect 5356 17060 5408 17066
rect 6012 17054 6132 17082
rect 5356 17002 5408 17008
rect 4871 16892 5179 16901
rect 4871 16890 4877 16892
rect 4933 16890 4957 16892
rect 5013 16890 5037 16892
rect 5093 16890 5117 16892
rect 5173 16890 5179 16892
rect 4933 16838 4935 16890
rect 5115 16838 5117 16890
rect 4871 16836 4877 16838
rect 4933 16836 4957 16838
rect 5013 16836 5037 16838
rect 5093 16836 5117 16838
rect 5173 16836 5179 16838
rect 4871 16827 5179 16836
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4080 16046 4108 16118
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 5092 15978 5120 16186
rect 5276 15978 5304 16458
rect 6104 16114 6132 17054
rect 6748 16998 6776 17546
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7024 16998 7052 17206
rect 7104 17128 7156 17134
rect 7102 17096 7104 17105
rect 7196 17128 7248 17134
rect 7156 17096 7158 17105
rect 7196 17070 7248 17076
rect 7102 17031 7158 17040
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6748 16114 6776 16934
rect 7024 16454 7052 16934
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7116 16182 7144 17031
rect 7208 16726 7236 17070
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7300 16522 7328 18294
rect 8036 18290 8064 19178
rect 8128 18766 8156 19790
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 8220 19378 8248 19722
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8496 18970 8524 19654
rect 8588 19378 8616 19926
rect 9692 19786 9720 20402
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 8792 19612 9100 19621
rect 8792 19610 8798 19612
rect 8854 19610 8878 19612
rect 8934 19610 8958 19612
rect 9014 19610 9038 19612
rect 9094 19610 9100 19612
rect 8854 19558 8856 19610
rect 9036 19558 9038 19610
rect 8792 19556 8798 19558
rect 8854 19556 8878 19558
rect 8934 19556 8958 19558
rect 9014 19556 9038 19558
rect 9094 19556 9100 19558
rect 8792 19547 9100 19556
rect 9036 19440 9088 19446
rect 9036 19382 9088 19388
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8116 18760 8168 18766
rect 8300 18760 8352 18766
rect 8116 18702 8168 18708
rect 8220 18720 8300 18748
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7576 17610 7604 18022
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 4871 15804 5179 15813
rect 4871 15802 4877 15804
rect 4933 15802 4957 15804
rect 5013 15802 5037 15804
rect 5093 15802 5117 15804
rect 5173 15802 5179 15804
rect 4933 15750 4935 15802
rect 5115 15750 5117 15802
rect 4871 15748 4877 15750
rect 4933 15748 4957 15750
rect 5013 15748 5037 15750
rect 5093 15748 5117 15750
rect 5173 15748 5179 15750
rect 4871 15739 5179 15748
rect 6104 15706 6132 16050
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3712 14006 3740 14214
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3068 13110 3188 13138
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2884 11150 2912 11766
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 9722 2360 10610
rect 2608 10606 2636 10950
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2700 10266 2728 10474
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2884 10146 2912 11086
rect 3068 10266 3096 13110
rect 3252 12850 3280 13126
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3160 12442 3188 12650
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3160 12306 3188 12378
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3252 12170 3280 12650
rect 3344 12374 3372 13194
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12850 3464 13126
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3252 11762 3280 12106
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10810 3464 10950
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10520 3188 10610
rect 3424 10532 3476 10538
rect 3160 10492 3424 10520
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2792 10118 2912 10146
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2792 9586 2820 10118
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2228 9580 2280 9586
rect 2780 9580 2832 9586
rect 2228 9522 2280 9528
rect 2700 9540 2780 9568
rect 2240 8974 2268 9522
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2056 8498 2084 8910
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2700 6798 2728 9540
rect 2780 9522 2832 9528
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2792 8498 2820 8910
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2792 8090 2820 8434
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 7886 2912 9930
rect 3068 9586 3096 10202
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 8838 3004 9318
rect 3068 9042 3096 9386
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9110 3188 9318
rect 3252 9110 3280 10492
rect 3424 10474 3476 10480
rect 3528 10266 3556 13874
rect 3712 12850 3740 13942
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3712 12646 3740 12786
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3988 12238 4016 12922
rect 4080 12918 4108 15506
rect 6748 15314 6776 16050
rect 6748 15286 6960 15314
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4448 13870 4476 14214
rect 4540 13938 4568 14758
rect 4871 14716 5179 14725
rect 4871 14714 4877 14716
rect 4933 14714 4957 14716
rect 5013 14714 5037 14716
rect 5093 14714 5117 14716
rect 5173 14714 5179 14716
rect 4933 14662 4935 14714
rect 5115 14662 5117 14714
rect 4871 14660 4877 14662
rect 4933 14660 4957 14662
rect 5013 14660 5037 14662
rect 5093 14660 5117 14662
rect 5173 14660 5179 14662
rect 4871 14651 5179 14660
rect 5644 14006 5672 14826
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4264 13394 4292 13806
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 4871 13628 5179 13637
rect 4871 13626 4877 13628
rect 4933 13626 4957 13628
rect 5013 13626 5037 13628
rect 5093 13626 5117 13628
rect 5173 13626 5179 13628
rect 4933 13574 4935 13626
rect 5115 13574 5117 13626
rect 4871 13572 4877 13574
rect 4933 13572 4957 13574
rect 5013 13572 5037 13574
rect 5093 13572 5117 13574
rect 5173 13572 5179 13574
rect 4871 13563 5179 13572
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 5368 13326 5396 13670
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 4068 12912 4120 12918
rect 4436 12912 4488 12918
rect 4120 12872 4200 12900
rect 4068 12854 4120 12860
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4080 11898 4108 12174
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2976 8362 3004 8774
rect 3068 8634 3096 8774
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7410 2912 7686
rect 2976 7546 3004 8298
rect 3252 7886 3280 8910
rect 3344 8906 3372 9998
rect 3528 9110 3556 10202
rect 3620 10062 3648 11698
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10810 4016 11086
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4172 10198 4200 12872
rect 4436 12854 4488 12860
rect 4448 11694 4476 12854
rect 4871 12540 5179 12549
rect 4871 12538 4877 12540
rect 4933 12538 4957 12540
rect 5013 12538 5037 12540
rect 5093 12538 5117 12540
rect 5173 12538 5179 12540
rect 4933 12486 4935 12538
rect 5115 12486 5117 12538
rect 4871 12484 4877 12486
rect 4933 12484 4957 12486
rect 5013 12484 5037 12486
rect 5093 12484 5117 12486
rect 5173 12484 5179 12486
rect 4871 12475 5179 12484
rect 5552 12306 5580 13126
rect 5828 12986 5856 13126
rect 5920 12986 5948 13466
rect 6012 13394 6040 13670
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12442 5672 12786
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3712 8974 3740 9522
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 8498 3372 8842
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 3068 6934 3096 7482
rect 3344 7426 3372 8434
rect 3804 8362 3832 10134
rect 4632 10062 4660 11630
rect 4724 11354 4752 11698
rect 5736 11694 5764 12718
rect 6104 12434 6132 14894
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6380 12442 6408 14486
rect 6656 14414 6684 14894
rect 6932 14890 6960 15286
rect 7116 15026 7144 16118
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14006 6776 14214
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6748 13802 6776 13942
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12850 6500 13262
rect 6564 12918 6592 13670
rect 7116 13530 7144 14350
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6012 12406 6132 12434
rect 6368 12436 6420 12442
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 6012 11558 6040 12406
rect 6368 12378 6420 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 12170 6408 12242
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 4871 11452 5179 11461
rect 4871 11450 4877 11452
rect 4933 11450 4957 11452
rect 5013 11450 5037 11452
rect 5093 11450 5117 11452
rect 5173 11450 5179 11452
rect 4933 11398 4935 11450
rect 5115 11398 5117 11450
rect 4871 11396 4877 11398
rect 4933 11396 4957 11398
rect 5013 11396 5037 11398
rect 5093 11396 5117 11398
rect 5173 11396 5179 11398
rect 4871 11387 5179 11396
rect 6012 11354 6040 11494
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 4871 10364 5179 10373
rect 4871 10362 4877 10364
rect 4933 10362 4957 10364
rect 5013 10362 5037 10364
rect 5093 10362 5117 10364
rect 5173 10362 5179 10364
rect 4933 10310 4935 10362
rect 5115 10310 5117 10362
rect 4871 10308 4877 10310
rect 4933 10308 4957 10310
rect 5013 10308 5037 10310
rect 5093 10308 5117 10310
rect 5173 10308 5179 10310
rect 4871 10299 5179 10308
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 3896 8430 3924 9998
rect 5276 9994 5304 10406
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4172 9178 4200 9522
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4724 8974 4752 9318
rect 4871 9276 5179 9285
rect 4871 9274 4877 9276
rect 4933 9274 4957 9276
rect 5013 9274 5037 9276
rect 5093 9274 5117 9276
rect 5173 9274 5179 9276
rect 4933 9222 4935 9274
rect 5115 9222 5117 9274
rect 4871 9220 4877 9222
rect 4933 9220 4957 9222
rect 5013 9220 5037 9222
rect 5093 9220 5117 9222
rect 5173 9220 5179 9222
rect 4871 9211 5179 9220
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 5644 8906 5672 11154
rect 6012 11150 6040 11290
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 9178 5764 10610
rect 5828 9586 5856 11018
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 4632 8566 4660 8842
rect 5460 8634 5488 8842
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3252 7398 3372 7426
rect 3252 7342 3280 7398
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 3344 6798 3372 7210
rect 3804 6866 3832 8298
rect 3896 7750 3924 8366
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 6322 4016 6734
rect 4172 6458 4200 7278
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4264 7002 4292 7210
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4356 6390 4384 6734
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4448 6322 4476 7142
rect 4632 6458 4660 8502
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5724 8492 5776 8498
rect 5828 8480 5856 9522
rect 5920 9518 5948 11018
rect 6104 10266 6132 11018
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5920 8945 5948 9454
rect 5906 8936 5962 8945
rect 5906 8871 5962 8880
rect 6012 8498 6040 9862
rect 6104 9722 6132 10202
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6380 8498 6408 9590
rect 6472 9178 6500 10610
rect 6564 10062 6592 12718
rect 6656 12170 6684 13126
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6748 11762 6776 13262
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 11286 6684 11494
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9722 6592 9998
rect 6748 9926 6776 11698
rect 6840 11082 6868 13194
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12442 7052 12786
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 9994 6868 10406
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 5776 8452 5856 8480
rect 6000 8492 6052 8498
rect 5724 8434 5776 8440
rect 6000 8434 6052 8440
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 4871 8188 5179 8197
rect 4871 8186 4877 8188
rect 4933 8186 4957 8188
rect 5013 8186 5037 8188
rect 5093 8186 5117 8188
rect 5173 8186 5179 8188
rect 4933 8134 4935 8186
rect 5115 8134 5117 8186
rect 4871 8132 4877 8134
rect 4933 8132 4957 8134
rect 5013 8132 5037 8134
rect 5093 8132 5117 8134
rect 5173 8132 5179 8134
rect 4871 8123 5179 8132
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4871 7100 5179 7109
rect 4871 7098 4877 7100
rect 4933 7098 4957 7100
rect 5013 7098 5037 7100
rect 5093 7098 5117 7100
rect 5173 7098 5179 7100
rect 4933 7046 4935 7098
rect 5115 7046 5117 7098
rect 4871 7044 4877 7046
rect 4933 7044 4957 7046
rect 5013 7044 5037 7046
rect 5093 7044 5117 7046
rect 5173 7044 5179 7046
rect 4871 7035 5179 7044
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 5000 6322 5028 6802
rect 5276 6798 5304 7686
rect 5552 7342 5580 8366
rect 5644 7546 5672 8434
rect 5736 8294 5764 8434
rect 6656 8294 6684 8842
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5736 7410 5764 8230
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5368 7002 5396 7278
rect 5552 7002 5580 7278
rect 6380 7002 6408 7754
rect 6656 7478 6684 8230
rect 6932 7954 6960 9522
rect 7024 8090 7052 9522
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7116 7886 7144 8298
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6748 7410 6776 7686
rect 7024 7546 7052 7754
rect 7208 7750 7236 11018
rect 7300 9042 7328 16458
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15570 7512 15846
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7668 14482 7696 18158
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 8036 17814 8064 18022
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7746 17640 7802 17649
rect 7746 17575 7748 17584
rect 7800 17575 7802 17584
rect 7748 17546 7800 17552
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7656 14340 7708 14346
rect 7760 14328 7788 17546
rect 8128 17134 8156 18702
rect 8220 17338 8248 18720
rect 8300 18702 8352 18708
rect 8496 18426 8524 18906
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8312 17542 8340 17750
rect 8404 17678 8432 18294
rect 8588 18154 8616 19314
rect 9048 19174 9076 19382
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8680 18970 8708 19110
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8680 18154 8708 18634
rect 8792 18524 9100 18533
rect 8792 18522 8798 18524
rect 8854 18522 8878 18524
rect 8934 18522 8958 18524
rect 9014 18522 9038 18524
rect 9094 18522 9100 18524
rect 8854 18470 8856 18522
rect 9036 18470 9038 18522
rect 8792 18468 8798 18470
rect 8854 18468 8878 18470
rect 8934 18468 8958 18470
rect 9014 18468 9038 18470
rect 9094 18468 9100 18470
rect 8792 18459 9100 18468
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8588 18034 8616 18090
rect 8588 18006 8708 18034
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8128 16794 8156 17070
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8128 15910 8156 16730
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8220 15502 8248 16594
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8404 16046 8432 16186
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14414 8156 14758
rect 8312 14618 8340 15982
rect 8404 15706 8432 15982
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8404 14618 8432 15370
rect 8496 15026 8524 15914
rect 8588 15706 8616 17614
rect 8680 17082 8708 18006
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8792 17436 9100 17445
rect 8792 17434 8798 17436
rect 8854 17434 8878 17436
rect 8934 17434 8958 17436
rect 9014 17434 9038 17436
rect 9094 17434 9100 17436
rect 8854 17382 8856 17434
rect 9036 17382 9038 17434
rect 8792 17380 8798 17382
rect 8854 17380 8878 17382
rect 8934 17380 8958 17382
rect 9014 17380 9038 17382
rect 9094 17380 9100 17382
rect 8792 17371 9100 17380
rect 9140 17270 9168 17478
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 8680 17054 9168 17082
rect 8792 16348 9100 16357
rect 8792 16346 8798 16348
rect 8854 16346 8878 16348
rect 8934 16346 8958 16348
rect 9014 16346 9038 16348
rect 9094 16346 9100 16348
rect 8854 16294 8856 16346
rect 9036 16294 9038 16346
rect 8792 16292 8798 16294
rect 8854 16292 8878 16294
rect 8934 16292 8958 16294
rect 9014 16292 9038 16294
rect 9094 16292 9100 16294
rect 8792 16283 9100 16292
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8588 15162 8616 15370
rect 8792 15260 9100 15269
rect 8792 15258 8798 15260
rect 8854 15258 8878 15260
rect 8934 15258 8958 15260
rect 9014 15258 9038 15260
rect 9094 15258 9100 15260
rect 8854 15206 8856 15258
rect 9036 15206 9038 15258
rect 8792 15204 8798 15206
rect 8854 15204 8878 15206
rect 8934 15204 8958 15206
rect 9014 15204 9038 15206
rect 9094 15204 9100 15206
rect 8792 15195 9100 15204
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8680 14929 8708 14962
rect 8666 14920 8722 14929
rect 8666 14855 8722 14864
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7708 14300 7788 14328
rect 7656 14282 7708 14288
rect 7760 14006 7788 14300
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8128 13530 8156 13670
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7392 12646 7420 13262
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 11762 7420 12582
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7576 11150 7604 13262
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7760 11558 7788 11766
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7576 9382 7604 11086
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 9110 7604 9318
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8566 7328 8978
rect 7576 8922 7604 9046
rect 7576 8906 7696 8922
rect 7576 8900 7708 8906
rect 7576 8894 7656 8900
rect 7656 8842 7708 8848
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6564 6798 6592 7142
rect 6748 6798 6776 7346
rect 7668 6866 7696 8434
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7760 6798 7788 11494
rect 8128 11150 8156 13466
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8312 8974 8340 14418
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 9994 8616 10950
rect 8680 10538 8708 14855
rect 8792 14172 9100 14181
rect 8792 14170 8798 14172
rect 8854 14170 8878 14172
rect 8934 14170 8958 14172
rect 9014 14170 9038 14172
rect 9094 14170 9100 14172
rect 8854 14118 8856 14170
rect 9036 14118 9038 14170
rect 8792 14116 8798 14118
rect 8854 14116 8878 14118
rect 8934 14116 8958 14118
rect 9014 14116 9038 14118
rect 9094 14116 9100 14118
rect 8792 14107 9100 14116
rect 8792 13084 9100 13093
rect 8792 13082 8798 13084
rect 8854 13082 8878 13084
rect 8934 13082 8958 13084
rect 9014 13082 9038 13084
rect 9094 13082 9100 13084
rect 8854 13030 8856 13082
rect 9036 13030 9038 13082
rect 8792 13028 8798 13030
rect 8854 13028 8878 13030
rect 8934 13028 8958 13030
rect 9014 13028 9038 13030
rect 9094 13028 9100 13030
rect 8792 13019 9100 13028
rect 9140 12238 9168 17054
rect 9232 16114 9260 19382
rect 9324 18766 9352 19654
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9416 18630 9444 19110
rect 9508 18970 9536 19382
rect 9600 19378 9628 19654
rect 9692 19514 9720 19722
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9968 19378 9996 20266
rect 10060 19446 10088 20402
rect 10152 20398 10180 20810
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9496 18760 9548 18766
rect 9600 18748 9628 19178
rect 9548 18720 9628 18748
rect 9680 18760 9732 18766
rect 9496 18702 9548 18708
rect 9680 18702 9732 18708
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 18426 9444 18566
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9324 16726 9352 17614
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16726 9444 16934
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9232 16017 9260 16050
rect 9218 16008 9274 16017
rect 9218 15943 9274 15952
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9232 13938 9260 15846
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 13938 9352 14758
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12986 9352 13126
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8792 11996 9100 12005
rect 8792 11994 8798 11996
rect 8854 11994 8878 11996
rect 8934 11994 8958 11996
rect 9014 11994 9038 11996
rect 9094 11994 9100 11996
rect 8854 11942 8856 11994
rect 9036 11942 9038 11994
rect 8792 11940 8798 11942
rect 8854 11940 8878 11942
rect 8934 11940 8958 11942
rect 9014 11940 9038 11942
rect 9094 11940 9100 11942
rect 8792 11931 9100 11940
rect 8792 10908 9100 10917
rect 8792 10906 8798 10908
rect 8854 10906 8878 10908
rect 8934 10906 8958 10908
rect 9014 10906 9038 10908
rect 9094 10906 9100 10908
rect 8854 10854 8856 10906
rect 9036 10854 9038 10906
rect 8792 10852 8798 10854
rect 8854 10852 8878 10854
rect 8934 10852 8958 10854
rect 9014 10852 9038 10854
rect 9094 10852 9100 10854
rect 8792 10843 9100 10852
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8792 9820 9100 9829
rect 8792 9818 8798 9820
rect 8854 9818 8878 9820
rect 8934 9818 8958 9820
rect 9014 9818 9038 9820
rect 9094 9818 9100 9820
rect 8854 9766 8856 9818
rect 9036 9766 9038 9818
rect 8792 9764 8798 9766
rect 8854 9764 8878 9766
rect 8934 9764 8958 9766
rect 9014 9764 9038 9766
rect 9094 9764 9100 9766
rect 8792 9755 9100 9764
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 8300 8968 8352 8974
rect 8484 8968 8536 8974
rect 8300 8910 8352 8916
rect 8404 8928 8484 8956
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7944 8498 7972 8774
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8128 7274 8156 8774
rect 8312 8090 8340 8910
rect 8404 8634 8432 8928
rect 8484 8910 8536 8916
rect 8792 8732 9100 8741
rect 8792 8730 8798 8732
rect 8854 8730 8878 8732
rect 8934 8730 8958 8732
rect 9014 8730 9038 8732
rect 9094 8730 9100 8732
rect 8854 8678 8856 8730
rect 9036 8678 9038 8730
rect 8792 8676 8798 8678
rect 8854 8676 8878 8678
rect 8934 8676 8958 8678
rect 9014 8676 9038 8678
rect 9094 8676 9100 8678
rect 8792 8667 9100 8676
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8312 7410 8340 8026
rect 8404 7410 8432 8570
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8496 8412 8524 8502
rect 8760 8424 8812 8430
rect 8496 8384 8760 8412
rect 8760 8366 8812 8372
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 7478 8708 7686
rect 8792 7644 9100 7653
rect 8792 7642 8798 7644
rect 8854 7642 8878 7644
rect 8934 7642 8958 7644
rect 9014 7642 9038 7644
rect 9094 7642 9100 7644
rect 8854 7590 8856 7642
rect 9036 7590 9038 7642
rect 8792 7588 8798 7590
rect 8854 7588 8878 7590
rect 8934 7588 8958 7590
rect 9014 7588 9038 7590
rect 9094 7588 9100 7590
rect 8792 7579 9100 7588
rect 9140 7546 9168 9046
rect 9324 7732 9352 9590
rect 9416 8974 9444 13194
rect 9508 12832 9536 18702
rect 9692 18290 9720 18702
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18358 9996 18566
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 10060 18086 10088 19382
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17882 10088 18022
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10244 17814 10272 20266
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10428 18766 10456 19314
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10428 18426 10456 18702
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10612 17814 10640 18770
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9692 17066 9720 17206
rect 9784 17134 9812 17478
rect 9876 17338 9904 17614
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9968 17270 9996 17614
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9876 17082 9904 17138
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9692 16658 9720 17002
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9680 16448 9732 16454
rect 9784 16436 9812 17070
rect 9876 17054 9996 17082
rect 9968 16590 9996 17054
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16794 10088 16934
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9732 16408 9812 16436
rect 9680 16390 9732 16396
rect 9588 16176 9640 16182
rect 9586 16144 9588 16153
rect 9640 16144 9642 16153
rect 9586 16079 9642 16088
rect 10152 15502 10180 17206
rect 10244 16658 10272 17750
rect 10414 16688 10470 16697
rect 10232 16652 10284 16658
rect 10284 16612 10364 16640
rect 10414 16623 10416 16632
rect 10232 16594 10284 16600
rect 10336 16182 10364 16612
rect 10468 16623 10470 16632
rect 10416 16594 10468 16600
rect 10428 16522 10456 16594
rect 10796 16590 10824 20334
rect 10980 19718 11008 20402
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10888 18970 10916 19314
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 11072 18902 11100 21247
rect 11716 20534 11744 21247
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19446 11192 19654
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11150 18728 11206 18737
rect 11072 18290 11100 18702
rect 11150 18663 11152 18672
rect 11204 18663 11206 18672
rect 11152 18634 11204 18640
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11164 17814 11192 18226
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11164 17678 11192 17750
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 11072 17241 11100 17546
rect 11256 17270 11284 19790
rect 11808 19718 11836 21383
rect 13082 21176 13138 21185
rect 13082 21111 13138 21120
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 17678 11376 18566
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11440 17882 11468 18226
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11244 17264 11296 17270
rect 11058 17232 11114 17241
rect 11244 17206 11296 17212
rect 11058 17167 11060 17176
rect 11112 17167 11114 17176
rect 11060 17138 11112 17144
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 10980 16250 11008 16934
rect 11440 16658 11468 17818
rect 11716 17814 11744 18022
rect 11704 17808 11756 17814
rect 11702 17776 11704 17785
rect 11756 17776 11758 17785
rect 11702 17711 11758 17720
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11808 16998 11836 17206
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 14414 9628 14758
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9692 14278 9720 14962
rect 9968 14618 9996 15030
rect 10152 14890 10180 15438
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9784 14414 9812 14486
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 14074 9720 14214
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 10152 13530 10180 14826
rect 10520 14822 10548 15846
rect 10612 15366 10640 15914
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 10704 15638 10732 15846
rect 11348 15706 11376 15846
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 11256 15570 11284 15642
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10520 13530 10548 14010
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9588 12844 9640 12850
rect 9508 12804 9588 12832
rect 9588 12786 9640 12792
rect 9600 12322 9628 12786
rect 9692 12442 9720 13262
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9600 12294 9720 12322
rect 9692 11150 9720 12294
rect 9784 11354 9812 13262
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 11150 9904 12786
rect 10612 12782 10640 15302
rect 11440 15094 11468 16390
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11532 15570 11560 15982
rect 11624 15638 11652 16526
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15434 11560 15506
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11716 15026 11744 16050
rect 11808 15910 11836 16934
rect 11900 16590 11928 18838
rect 11992 17882 12020 20402
rect 12176 19854 12204 20402
rect 12713 20156 13021 20165
rect 12713 20154 12719 20156
rect 12775 20154 12799 20156
rect 12855 20154 12879 20156
rect 12935 20154 12959 20156
rect 13015 20154 13021 20156
rect 12775 20102 12777 20154
rect 12957 20102 12959 20154
rect 12713 20100 12719 20102
rect 12775 20100 12799 20102
rect 12855 20100 12879 20102
rect 12935 20100 12959 20102
rect 13015 20100 13021 20102
rect 12713 20091 13021 20100
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 12084 19378 12112 19722
rect 12176 19514 12204 19790
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11992 16114 12020 17478
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 12084 16046 12112 19314
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12360 18193 12388 18226
rect 12346 18184 12402 18193
rect 12346 18119 12402 18128
rect 12452 18086 12480 18566
rect 12544 18290 12572 18702
rect 12636 18426 12664 19790
rect 13096 19446 13124 21111
rect 13542 20632 13598 20641
rect 13542 20567 13544 20576
rect 13596 20567 13598 20576
rect 13544 20538 13596 20544
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 12713 19068 13021 19077
rect 12713 19066 12719 19068
rect 12775 19066 12799 19068
rect 12855 19066 12879 19068
rect 12935 19066 12959 19068
rect 13015 19066 13021 19068
rect 12775 19014 12777 19066
rect 12957 19014 12959 19066
rect 12713 19012 12719 19014
rect 12775 19012 12799 19014
rect 12855 19012 12879 19014
rect 12935 19012 12959 19014
rect 13015 19012 13021 19014
rect 12713 19003 13021 19012
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12728 18170 12756 18566
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12544 18142 12756 18170
rect 12912 18154 12940 18226
rect 12900 18148 12952 18154
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12544 17610 12572 18142
rect 12900 18090 12952 18096
rect 12713 17980 13021 17989
rect 12713 17978 12719 17980
rect 12775 17978 12799 17980
rect 12855 17978 12879 17980
rect 12935 17978 12959 17980
rect 13015 17978 13021 17980
rect 12775 17926 12777 17978
rect 12957 17926 12959 17978
rect 12713 17924 12719 17926
rect 12775 17924 12799 17926
rect 12855 17924 12879 17926
rect 12935 17924 12959 17926
rect 13015 17924 13021 17926
rect 12713 17915 13021 17924
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12728 17678 12756 17750
rect 12716 17672 12768 17678
rect 12636 17632 12716 17660
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12176 16046 12204 17002
rect 12268 16590 12296 17138
rect 12452 16794 12480 17546
rect 12544 17338 12572 17546
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11900 14890 11928 15438
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10704 13938 10732 14758
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10796 13258 10824 14554
rect 11900 14482 11928 14826
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 11440 13190 11468 14282
rect 11624 14074 11652 14282
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11518 13424 11574 13433
rect 11518 13359 11574 13368
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 10062 9720 10406
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9678 9616 9734 9625
rect 9678 9551 9680 9560
rect 9732 9551 9734 9560
rect 9680 9522 9732 9528
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7744 9456 7750
rect 9324 7704 9404 7732
rect 9404 7686 9456 7692
rect 9508 7546 9536 8026
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9600 7478 9628 7686
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8312 7290 8340 7346
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8220 7262 8340 7290
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 5276 6390 5304 6734
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 8128 6254 8156 7210
rect 8220 6798 8248 7262
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8404 6338 8432 7346
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 6866 8616 7142
rect 9416 6866 9444 7414
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 8792 6556 9100 6565
rect 8792 6554 8798 6556
rect 8854 6554 8878 6556
rect 8934 6554 8958 6556
rect 9014 6554 9038 6556
rect 9094 6554 9100 6556
rect 8854 6502 8856 6554
rect 9036 6502 9038 6554
rect 8792 6500 8798 6502
rect 8854 6500 8878 6502
rect 8934 6500 8958 6502
rect 9014 6500 9038 6502
rect 9094 6500 9100 6502
rect 8792 6491 9100 6500
rect 8312 6322 8616 6338
rect 9508 6322 9536 6734
rect 9600 6662 9628 7278
rect 9692 6866 9720 8842
rect 9784 8430 9812 10542
rect 9876 9110 9904 11086
rect 9968 9518 9996 12242
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10060 10810 10088 11018
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10152 10266 10180 11630
rect 10244 11150 10272 12582
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 11354 10456 12106
rect 11164 11762 11192 12174
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10140 10260 10192 10266
rect 10060 10220 10140 10248
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9968 8498 9996 9454
rect 10060 8838 10088 10220
rect 10140 10202 10192 10208
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10152 8537 10180 9522
rect 10244 9178 10272 10610
rect 10414 9616 10470 9625
rect 10324 9580 10376 9586
rect 10414 9551 10416 9560
rect 10324 9522 10376 9528
rect 10468 9551 10470 9560
rect 10416 9522 10468 9528
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8566 10272 8774
rect 10336 8634 10364 9522
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10888 8566 10916 9046
rect 10232 8560 10284 8566
rect 10138 8528 10194 8537
rect 9956 8492 10008 8498
rect 10232 8502 10284 8508
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10138 8463 10194 8472
rect 9956 8434 10008 8440
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9784 6662 9812 7346
rect 9968 7274 9996 7822
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7478 10180 7754
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 10152 6458 10180 7414
rect 10244 6798 10272 7958
rect 10336 7410 10364 8230
rect 10980 7478 11008 8230
rect 11072 7886 11100 11086
rect 11164 10062 11192 11698
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11348 9518 11376 9930
rect 11440 9625 11468 13126
rect 11532 12850 11560 13359
rect 11992 13326 12020 15030
rect 12084 14618 12112 15982
rect 12176 15502 12204 15982
rect 12268 15502 12296 16526
rect 12544 16250 12572 17138
rect 12636 16998 12664 17632
rect 12716 17614 12768 17620
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17338 12756 17478
rect 12912 17338 12940 17546
rect 13096 17513 13124 18634
rect 13188 17610 13216 19314
rect 13464 18902 13492 19314
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13268 18760 13320 18766
rect 13360 18760 13412 18766
rect 13268 18702 13320 18708
rect 13358 18728 13360 18737
rect 13412 18728 13414 18737
rect 13280 17610 13308 18702
rect 13358 18663 13414 18672
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 13082 17504 13138 17513
rect 13082 17439 13138 17448
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12713 16892 13021 16901
rect 12713 16890 12719 16892
rect 12775 16890 12799 16892
rect 12855 16890 12879 16892
rect 12935 16890 12959 16892
rect 13015 16890 13021 16892
rect 12775 16838 12777 16890
rect 12957 16838 12959 16890
rect 12713 16836 12719 16838
rect 12775 16836 12799 16838
rect 12855 16836 12879 16838
rect 12935 16836 12959 16838
rect 13015 16836 13021 16838
rect 12713 16827 13021 16836
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12636 15570 12664 16662
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13004 15978 13032 16526
rect 13096 16454 13124 17439
rect 13280 17218 13308 17546
rect 13188 17190 13308 17218
rect 13372 17202 13400 18663
rect 13464 17678 13492 18838
rect 13556 18766 13584 19654
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13648 18426 13676 20402
rect 13832 20330 13860 21383
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 14200 20058 14228 21383
rect 15856 20806 15884 21383
rect 27342 21040 27398 21049
rect 27342 20975 27398 20984
rect 17130 20904 17186 20913
rect 17130 20839 17186 20848
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 16634 20700 16942 20709
rect 16634 20698 16640 20700
rect 16696 20698 16720 20700
rect 16776 20698 16800 20700
rect 16856 20698 16880 20700
rect 16936 20698 16942 20700
rect 16696 20646 16698 20698
rect 16878 20646 16880 20698
rect 16634 20644 16640 20646
rect 16696 20644 16720 20646
rect 16776 20644 16800 20646
rect 16856 20644 16880 20646
rect 16936 20644 16942 20646
rect 16118 20632 16174 20641
rect 16634 20635 16942 20644
rect 16118 20567 16120 20576
rect 16172 20567 16174 20576
rect 17038 20632 17094 20641
rect 17038 20567 17040 20576
rect 16120 20538 16172 20544
rect 17092 20567 17094 20576
rect 17040 20538 17092 20544
rect 15384 20528 15436 20534
rect 15436 20476 15516 20482
rect 15384 20470 15516 20476
rect 15396 20454 15516 20470
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 13740 19417 13768 19790
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 13726 19408 13782 19417
rect 14660 19378 14688 19722
rect 13726 19343 13782 19352
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14476 18630 14504 19178
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18970 14596 19110
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14186 18184 14242 18193
rect 14186 18119 14242 18128
rect 14200 18086 14228 18119
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13740 17610 13768 18022
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13360 17196 13412 17202
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13082 16144 13138 16153
rect 13082 16079 13084 16088
rect 13136 16079 13138 16088
rect 13084 16050 13136 16056
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 12713 15804 13021 15813
rect 12713 15802 12719 15804
rect 12775 15802 12799 15804
rect 12855 15802 12879 15804
rect 12935 15802 12959 15804
rect 13015 15802 13021 15804
rect 12775 15750 12777 15802
rect 12957 15750 12959 15802
rect 12713 15748 12719 15750
rect 12775 15748 12799 15750
rect 12855 15748 12879 15750
rect 12935 15748 12959 15750
rect 13015 15748 13021 15750
rect 12713 15739 13021 15748
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12452 14278 12480 14962
rect 12713 14716 13021 14725
rect 12713 14714 12719 14716
rect 12775 14714 12799 14716
rect 12855 14714 12879 14716
rect 12935 14714 12959 14716
rect 13015 14714 13021 14716
rect 12775 14662 12777 14714
rect 12957 14662 12959 14714
rect 12713 14660 12719 14662
rect 12775 14660 12799 14662
rect 12855 14660 12879 14662
rect 12935 14660 12959 14662
rect 13015 14660 13021 14662
rect 12713 14651 13021 14660
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12728 14521 12756 14554
rect 12714 14512 12770 14521
rect 12714 14447 12770 14456
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12728 14074 12756 14282
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 13096 13977 13124 16050
rect 13188 15910 13216 17190
rect 13360 17138 13412 17144
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13372 16658 13400 17138
rect 13464 16726 13492 17138
rect 13648 17066 13676 17138
rect 13740 17066 13768 17546
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13188 14414 13216 15846
rect 13372 15434 13400 16118
rect 13464 16114 13492 16526
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13082 13968 13138 13977
rect 13082 13903 13138 13912
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13530 12664 13670
rect 12713 13628 13021 13637
rect 12713 13626 12719 13628
rect 12775 13626 12799 13628
rect 12855 13626 12879 13628
rect 12935 13626 12959 13628
rect 13015 13626 13021 13628
rect 12775 13574 12777 13626
rect 12957 13574 12959 13626
rect 12713 13572 12719 13574
rect 12775 13572 12799 13574
rect 12855 13572 12879 13574
rect 12935 13572 12959 13574
rect 13015 13572 13021 13574
rect 12713 13563 13021 13572
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12442 11560 12786
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 12084 12238 12112 13126
rect 12176 12918 12204 13262
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12713 12540 13021 12549
rect 12713 12538 12719 12540
rect 12775 12538 12799 12540
rect 12855 12538 12879 12540
rect 12935 12538 12959 12540
rect 13015 12538 13021 12540
rect 12775 12486 12777 12538
rect 12957 12486 12959 12538
rect 12713 12484 12719 12486
rect 12775 12484 12799 12486
rect 12855 12484 12879 12486
rect 12935 12484 12959 12486
rect 13015 12484 13021 12486
rect 12713 12475 13021 12484
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12452 11558 12480 12038
rect 12544 11830 12572 12038
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11900 10674 11928 11086
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11888 10668 11940 10674
rect 11940 10628 12020 10656
rect 11888 10610 11940 10616
rect 11426 9616 11482 9625
rect 11426 9551 11482 9560
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 8566 11652 9318
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11716 8362 11744 10610
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 8974 11836 10406
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11900 9586 11928 9862
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11992 9382 12020 10628
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 12452 8974 12480 11494
rect 12713 11452 13021 11461
rect 12713 11450 12719 11452
rect 12775 11450 12799 11452
rect 12855 11450 12879 11452
rect 12935 11450 12959 11452
rect 13015 11450 13021 11452
rect 12775 11398 12777 11450
rect 12957 11398 12959 11450
rect 12713 11396 12719 11398
rect 12775 11396 12799 11398
rect 12855 11396 12879 11398
rect 12935 11396 12959 11398
rect 13015 11396 13021 11398
rect 12713 11387 13021 11396
rect 13096 10742 13124 13903
rect 13372 13870 13400 14894
rect 13464 14618 13492 16050
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 15026 13584 15302
rect 13648 15026 13676 15438
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13726 15056 13782 15065
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13636 15020 13688 15026
rect 13924 15026 13952 15370
rect 13726 14991 13782 15000
rect 13912 15020 13964 15026
rect 13636 14962 13688 14968
rect 13740 14958 13768 14991
rect 13912 14962 13964 14968
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13648 14346 13676 14758
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 13870 13676 14282
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 13938 13860 14214
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 14108 13462 14136 14894
rect 14200 14482 14228 18022
rect 14292 17678 14320 18226
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14384 17814 14412 18022
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14554 17776 14610 17785
rect 14554 17711 14610 17720
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14384 15638 14412 16594
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14384 15026 14412 15574
rect 14476 15434 14504 17070
rect 14568 16794 14596 17711
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14660 16182 14688 19314
rect 14752 18834 14780 19790
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14752 18034 14780 18770
rect 15028 18766 15056 19994
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15304 19446 15332 19858
rect 15396 19854 15424 20334
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15488 18766 15516 20454
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 19786 15792 20198
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 18426 15516 18702
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14752 18006 14872 18034
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14752 17202 14780 17818
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14752 16794 14780 17138
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14844 16726 14872 18006
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14832 16584 14884 16590
rect 14830 16552 14832 16561
rect 14884 16552 14886 16561
rect 14830 16487 14886 16496
rect 14648 16176 14700 16182
rect 14648 16118 14700 16124
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14660 14890 14688 16118
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14660 14618 14688 14826
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14370 14512 14426 14521
rect 14188 14476 14240 14482
rect 14370 14447 14426 14456
rect 14188 14418 14240 14424
rect 14384 14414 14412 14447
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13174 13016 13230 13025
rect 13174 12951 13230 12960
rect 13188 12850 13216 12951
rect 13464 12850 13492 13126
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13556 12442 13584 12582
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13648 12238 13676 13126
rect 13740 12442 13768 13262
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12713 10364 13021 10373
rect 12713 10362 12719 10364
rect 12775 10362 12799 10364
rect 12855 10362 12879 10364
rect 12935 10362 12959 10364
rect 13015 10362 13021 10364
rect 12775 10310 12777 10362
rect 12957 10310 12959 10362
rect 12713 10308 12719 10310
rect 12775 10308 12799 10310
rect 12855 10308 12879 10310
rect 12935 10308 12959 10310
rect 13015 10308 13021 10310
rect 12713 10299 13021 10308
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 12544 9518 12572 9930
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9654 12940 9862
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 11796 8968 11848 8974
rect 11980 8968 12032 8974
rect 11796 8910 11848 8916
rect 11900 8928 11980 8956
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11348 7546 11376 7822
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 11624 7342 11652 8298
rect 11900 7886 11928 8928
rect 11980 8910 12032 8916
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12176 8498 12204 8842
rect 12360 8566 12388 8842
rect 12544 8634 12572 9454
rect 12636 9178 12664 9522
rect 12713 9276 13021 9285
rect 12713 9274 12719 9276
rect 12775 9274 12799 9276
rect 12855 9274 12879 9276
rect 12935 9274 12959 9276
rect 13015 9274 13021 9276
rect 12775 9222 12777 9274
rect 12957 9222 12959 9274
rect 12713 9220 12719 9222
rect 12775 9220 12799 9222
rect 12855 9220 12879 9222
rect 12935 9220 12959 9222
rect 13015 9220 13021 9222
rect 12713 9211 13021 9220
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12164 8492 12216 8498
rect 12216 8452 12296 8480
rect 12164 8434 12216 8440
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12268 7546 12296 8452
rect 12636 8430 12664 9114
rect 13096 9042 13124 9522
rect 13188 9178 13216 9930
rect 13280 9586 13308 11494
rect 13464 11098 13492 12106
rect 13924 12102 13952 12786
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14108 11762 14136 13398
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14280 12368 14332 12374
rect 14278 12336 14280 12345
rect 14332 12336 14334 12345
rect 14278 12271 14334 12280
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13648 11286 13676 11698
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 14384 11150 14412 13126
rect 14568 12918 14596 13330
rect 14660 13297 14688 13466
rect 14752 13326 14780 13670
rect 14740 13320 14792 13326
rect 14646 13288 14702 13297
rect 14740 13262 14792 13268
rect 14646 13223 14702 13232
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14476 12238 14504 12650
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14660 11830 14688 13223
rect 14738 13016 14794 13025
rect 14738 12951 14794 12960
rect 14648 11824 14700 11830
rect 14462 11792 14518 11801
rect 14648 11766 14700 11772
rect 14462 11727 14464 11736
rect 14516 11727 14518 11736
rect 14464 11698 14516 11704
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14372 11144 14424 11150
rect 13634 11112 13690 11121
rect 13464 11070 13634 11098
rect 14372 11086 14424 11092
rect 13634 11047 13690 11056
rect 13648 10538 13676 11047
rect 14568 11014 14596 11630
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 9625 13584 10406
rect 13740 9994 13768 10542
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13542 9616 13598 9625
rect 13268 9580 13320 9586
rect 13542 9551 13598 9560
rect 13268 9522 13320 9528
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 12728 8498 12756 8910
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12713 8188 13021 8197
rect 12713 8186 12719 8188
rect 12775 8186 12799 8188
rect 12855 8186 12879 8188
rect 12935 8186 12959 8188
rect 13015 8186 13021 8188
rect 12775 8134 12777 8186
rect 12957 8134 12959 8186
rect 12713 8132 12719 8134
rect 12775 8132 12799 8134
rect 12855 8132 12879 8134
rect 12935 8132 12959 8134
rect 13015 8132 13021 8134
rect 12713 8123 13021 8132
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 13188 7410 13216 7686
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6798 10456 7142
rect 12268 6866 12296 7346
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12713 7100 13021 7109
rect 12713 7098 12719 7100
rect 12775 7098 12799 7100
rect 12855 7098 12879 7100
rect 12935 7098 12959 7100
rect 13015 7098 13021 7100
rect 12775 7046 12777 7098
rect 12957 7046 12959 7098
rect 12713 7044 12719 7046
rect 12775 7044 12799 7046
rect 12855 7044 12879 7046
rect 12935 7044 12959 7046
rect 13015 7044 13021 7046
rect 12713 7035 13021 7044
rect 13096 7002 13124 7278
rect 13464 7274 13492 8570
rect 13556 7410 13584 9551
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13648 8945 13676 9046
rect 13634 8936 13690 8945
rect 13634 8871 13690 8880
rect 13740 7750 13768 9930
rect 14476 9654 14504 10678
rect 14568 9722 14596 10950
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14476 9042 14504 9590
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8566 14504 8978
rect 14660 8634 14688 11494
rect 14752 10742 14780 12951
rect 14844 12238 14872 14010
rect 14936 13734 14964 18226
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 15028 17921 15056 18090
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15014 17912 15070 17921
rect 15304 17882 15332 18022
rect 15014 17847 15070 17856
rect 15200 17876 15252 17882
rect 15028 16998 15056 17847
rect 15200 17818 15252 17824
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17513 15148 17614
rect 15106 17504 15162 17513
rect 15106 17439 15162 17448
rect 15016 16992 15068 16998
rect 15212 16969 15240 17818
rect 15396 17678 15424 18022
rect 15488 17921 15516 18158
rect 15474 17912 15530 17921
rect 15474 17847 15530 17856
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15016 16934 15068 16940
rect 15198 16960 15254 16969
rect 15198 16895 15254 16904
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15120 15706 15148 16594
rect 15108 15700 15160 15706
rect 15028 15660 15108 15688
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13326 14964 13670
rect 15028 13462 15056 15660
rect 15108 15642 15160 15648
rect 15212 15502 15240 16895
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 15028 12832 15056 13398
rect 15120 13190 15148 14962
rect 15212 13462 15240 15438
rect 15488 15366 15516 16050
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15396 14414 15424 14962
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 14006 15332 14214
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15396 13938 15424 14350
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15292 13864 15344 13870
rect 15488 13818 15516 15302
rect 15580 14074 15608 18634
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15672 18086 15700 18226
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15764 16794 15792 19722
rect 16408 19514 16436 20402
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16634 19612 16942 19621
rect 16634 19610 16640 19612
rect 16696 19610 16720 19612
rect 16776 19610 16800 19612
rect 16856 19610 16880 19612
rect 16936 19610 16942 19612
rect 16696 19558 16698 19610
rect 16878 19558 16880 19610
rect 16634 19556 16640 19558
rect 16696 19556 16720 19558
rect 16776 19556 16800 19558
rect 16856 19556 16880 19558
rect 16936 19556 16942 19558
rect 16634 19547 16942 19556
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 17052 19378 17080 19654
rect 17144 19514 17172 20839
rect 24476 20700 24784 20709
rect 24476 20698 24482 20700
rect 24538 20698 24562 20700
rect 24618 20698 24642 20700
rect 24698 20698 24722 20700
rect 24778 20698 24784 20700
rect 24538 20646 24540 20698
rect 24720 20646 24722 20698
rect 24476 20644 24482 20646
rect 24538 20644 24562 20646
rect 24618 20644 24642 20646
rect 24698 20644 24722 20646
rect 24778 20644 24784 20646
rect 24476 20635 24784 20644
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 17420 20330 17448 20470
rect 27356 20466 27384 20975
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17420 19854 17448 20266
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18766 15884 19110
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15844 18624 15896 18630
rect 15948 18612 15976 18702
rect 16500 18630 16528 19314
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 18766 17172 19110
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 15896 18584 15976 18612
rect 16304 18624 16356 18630
rect 15844 18566 15896 18572
rect 16304 18566 16356 18572
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 15856 18290 15884 18566
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15948 18086 15976 18226
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17134 16160 18022
rect 16210 17912 16266 17921
rect 16210 17847 16266 17856
rect 16224 17746 16252 17847
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16316 17678 16344 18566
rect 16634 18524 16942 18533
rect 16634 18522 16640 18524
rect 16696 18522 16720 18524
rect 16776 18522 16800 18524
rect 16856 18522 16880 18524
rect 16936 18522 16942 18524
rect 16696 18470 16698 18522
rect 16878 18470 16880 18522
rect 16634 18468 16640 18470
rect 16696 18468 16720 18470
rect 16776 18468 16800 18470
rect 16856 18468 16880 18470
rect 16936 18468 16942 18470
rect 16634 18459 16942 18468
rect 17420 18086 17448 18906
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17678 17448 18022
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 16500 17338 16528 17614
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 16634 17436 16942 17445
rect 16634 17434 16640 17436
rect 16696 17434 16720 17436
rect 16776 17434 16800 17436
rect 16856 17434 16880 17436
rect 16936 17434 16942 17436
rect 16696 17382 16698 17434
rect 16878 17382 16880 17434
rect 16634 17380 16640 17382
rect 16696 17380 16720 17382
rect 16776 17380 16800 17382
rect 16856 17380 16880 17382
rect 16936 17380 16942 17382
rect 16634 17371 16942 17380
rect 17144 17338 17172 17546
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16794 16068 16934
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16394 16688 16450 16697
rect 16394 16623 16450 16632
rect 16408 16590 16436 16623
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 15672 16250 15700 16526
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 14890 15792 15438
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15344 13812 15516 13818
rect 15292 13806 15516 13812
rect 15304 13790 15516 13806
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15108 12844 15160 12850
rect 15028 12804 15108 12832
rect 15108 12786 15160 12792
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15212 12374 15240 12650
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14844 11898 14872 12174
rect 15304 12170 15332 13670
rect 15396 13530 15424 13790
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15396 12442 15424 13466
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15488 13326 15516 13398
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15212 11830 15240 12106
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 8974 14780 9318
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14464 8560 14516 8566
rect 14186 8528 14242 8537
rect 14096 8492 14148 8498
rect 14464 8502 14516 8508
rect 14186 8463 14188 8472
rect 14096 8434 14148 8440
rect 14240 8463 14242 8472
rect 14188 8434 14240 8440
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7410 13860 7686
rect 14108 7546 14136 8434
rect 14476 7954 14504 8502
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14568 7886 14596 8298
rect 14660 8294 14688 8570
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 11532 6390 11560 6734
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11992 6322 12020 6598
rect 8300 6316 8628 6322
rect 8352 6310 8576 6316
rect 8300 6258 8352 6264
rect 8576 6258 8628 6264
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 4871 6012 5179 6021
rect 4871 6010 4877 6012
rect 4933 6010 4957 6012
rect 5013 6010 5037 6012
rect 5093 6010 5117 6012
rect 5173 6010 5179 6012
rect 4933 5958 4935 6010
rect 5115 5958 5117 6010
rect 4871 5956 4877 5958
rect 4933 5956 4957 5958
rect 5013 5956 5037 5958
rect 5093 5956 5117 5958
rect 5173 5956 5179 5958
rect 4871 5947 5179 5956
rect 11992 5914 12020 6258
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12176 5710 12204 6734
rect 12452 6662 12480 6802
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6118 12480 6598
rect 13740 6458 13768 7346
rect 13832 6934 13860 7346
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12713 6012 13021 6021
rect 12713 6010 12719 6012
rect 12775 6010 12799 6012
rect 12855 6010 12879 6012
rect 12935 6010 12959 6012
rect 13015 6010 13021 6012
rect 12775 5958 12777 6010
rect 12957 5958 12959 6010
rect 12713 5956 12719 5958
rect 12775 5956 12799 5958
rect 12855 5956 12879 5958
rect 12935 5956 12959 5958
rect 13015 5956 13021 5958
rect 12713 5947 13021 5956
rect 13188 5914 13216 6190
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13832 5846 13860 6870
rect 14844 6866 14872 11086
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 8634 14964 9998
rect 15028 9926 15056 10066
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15120 9466 15148 9930
rect 15212 9654 15240 11494
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15304 10810 15332 11290
rect 15396 11150 15424 12378
rect 15488 12306 15516 13262
rect 15580 13025 15608 13262
rect 15566 13016 15622 13025
rect 15672 12986 15700 13874
rect 15566 12951 15622 12960
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15764 12442 15792 14826
rect 15856 13734 15884 15982
rect 15948 14278 15976 16458
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 16132 15162 16160 16118
rect 16500 15910 16528 16526
rect 17512 16454 17540 20334
rect 18616 19786 18644 20402
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18604 19780 18656 19786
rect 18524 19740 18604 19768
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18426 18460 19110
rect 18524 18766 18552 19740
rect 18604 19722 18656 19728
rect 18602 19544 18658 19553
rect 18602 19479 18604 19488
rect 18656 19479 18658 19488
rect 18604 19450 18656 19456
rect 18708 19242 18736 19790
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18800 19378 18828 19654
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18708 18970 18736 19178
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18892 18834 18920 20198
rect 18984 20058 19012 20402
rect 20180 20058 20208 20402
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 19812 19910 20116 19938
rect 19812 19854 19840 19910
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19996 19718 20024 19790
rect 20088 19786 20116 19910
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18524 18426 18552 18702
rect 19536 18698 19564 19314
rect 20168 19304 20220 19310
rect 19614 19272 19670 19281
rect 20168 19246 20220 19252
rect 19614 19207 19670 19216
rect 19628 18902 19656 19207
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 18902 19748 19110
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19708 18896 19760 18902
rect 19708 18838 19760 18844
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 17105 17632 17614
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17202 17724 17478
rect 17788 17270 17816 17682
rect 18432 17678 18460 18362
rect 18788 18352 18840 18358
rect 18788 18294 18840 18300
rect 18800 18154 18828 18294
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 18800 17678 18828 18090
rect 18892 17678 18920 18566
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 19260 17610 19288 18158
rect 19536 18154 19564 18634
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19536 17882 19564 18090
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 17590 17096 17646 17105
rect 17590 17031 17646 17040
rect 17776 16992 17828 16998
rect 18524 16969 18552 17138
rect 17776 16934 17828 16940
rect 18510 16960 18566 16969
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 16634 16348 16942 16357
rect 16634 16346 16640 16348
rect 16696 16346 16720 16348
rect 16776 16346 16800 16348
rect 16856 16346 16880 16348
rect 16936 16346 16942 16348
rect 16696 16294 16698 16346
rect 16878 16294 16880 16346
rect 16634 16292 16640 16294
rect 16696 16292 16720 16294
rect 16776 16292 16800 16294
rect 16856 16292 16880 16294
rect 16936 16292 16942 16294
rect 16634 16283 16942 16292
rect 17788 16114 17816 16934
rect 18510 16895 18566 16904
rect 18786 16960 18842 16969
rect 18786 16895 18842 16904
rect 18418 16416 18474 16425
rect 18418 16351 18474 16360
rect 18432 16182 18460 16351
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16500 15706 16528 15846
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16500 15026 16528 15302
rect 16634 15260 16942 15269
rect 16634 15258 16640 15260
rect 16696 15258 16720 15260
rect 16776 15258 16800 15260
rect 16856 15258 16880 15260
rect 16936 15258 16942 15260
rect 16696 15206 16698 15258
rect 16878 15206 16880 15258
rect 16634 15204 16640 15206
rect 16696 15204 16720 15206
rect 16776 15204 16800 15206
rect 16856 15204 16880 15206
rect 16936 15204 16942 15206
rect 16634 15195 16942 15204
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16960 14822 16988 14962
rect 17052 14890 17080 16050
rect 17696 15706 18000 15722
rect 17684 15700 18000 15706
rect 17736 15694 18000 15700
rect 17684 15642 17736 15648
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16316 14414 16344 14758
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15948 12714 15976 14214
rect 16634 14172 16942 14181
rect 16634 14170 16640 14172
rect 16696 14170 16720 14172
rect 16776 14170 16800 14172
rect 16856 14170 16880 14172
rect 16936 14170 16942 14172
rect 16696 14118 16698 14170
rect 16878 14118 16880 14170
rect 16634 14116 16640 14118
rect 16696 14116 16720 14118
rect 16776 14116 16800 14118
rect 16856 14116 16880 14118
rect 16936 14116 16942 14118
rect 16634 14107 16942 14116
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16132 13258 16160 13942
rect 17052 13938 17080 14826
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16132 12918 16160 13194
rect 16634 13084 16942 13093
rect 16634 13082 16640 13084
rect 16696 13082 16720 13084
rect 16776 13082 16800 13084
rect 16856 13082 16880 13084
rect 16936 13082 16942 13084
rect 16696 13030 16698 13082
rect 16878 13030 16880 13082
rect 16634 13028 16640 13030
rect 16696 13028 16720 13030
rect 16776 13028 16800 13030
rect 16856 13028 16880 13030
rect 16936 13028 16942 13030
rect 16634 13019 16942 13028
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11898 15516 12038
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15580 11762 15608 12310
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15580 11150 15608 11698
rect 15764 11694 15792 12378
rect 15856 12102 15884 12378
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15304 10266 15332 10610
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15396 9518 15424 10610
rect 15488 9586 15516 11018
rect 15672 10810 15700 11154
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15764 10674 15792 10950
rect 15856 10810 15884 11766
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15948 11082 15976 11494
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15580 10062 15608 10202
rect 15672 10198 15700 10610
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15200 9512 15252 9518
rect 15120 9460 15200 9466
rect 15120 9454 15252 9460
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15120 9438 15240 9454
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15120 8498 15148 8910
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15396 7546 15424 7754
rect 15948 7750 15976 9454
rect 16040 9178 16068 12786
rect 16132 11626 16160 12854
rect 17144 12442 17172 14758
rect 17328 13938 17356 15302
rect 17788 15162 17816 15302
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17972 15026 18000 15694
rect 18432 15434 18460 16118
rect 18800 15960 18828 16895
rect 19260 16561 19288 17546
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 17134 19380 17478
rect 19444 17202 19472 17750
rect 19628 17626 19656 18362
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19720 17814 19748 18022
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19708 17672 19760 17678
rect 19628 17620 19708 17626
rect 19628 17614 19760 17620
rect 19628 17598 19748 17614
rect 19812 17338 19840 18838
rect 20180 18086 20208 19246
rect 20272 18970 20300 20402
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20456 20058 20484 20198
rect 20555 20156 20863 20165
rect 20555 20154 20561 20156
rect 20617 20154 20641 20156
rect 20697 20154 20721 20156
rect 20777 20154 20801 20156
rect 20857 20154 20863 20156
rect 20617 20102 20619 20154
rect 20799 20102 20801 20154
rect 20555 20100 20561 20102
rect 20617 20100 20641 20102
rect 20697 20100 20721 20102
rect 20777 20100 20801 20102
rect 20857 20100 20863 20102
rect 20555 20091 20863 20100
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20916 19718 20944 20402
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 20058 22140 20334
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 21008 19514 21036 19926
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20364 18698 20392 19314
rect 20456 18766 20484 19314
rect 20555 19068 20863 19077
rect 20555 19066 20561 19068
rect 20617 19066 20641 19068
rect 20697 19066 20721 19068
rect 20777 19066 20801 19068
rect 20857 19066 20863 19068
rect 20617 19014 20619 19066
rect 20799 19014 20801 19066
rect 20555 19012 20561 19014
rect 20617 19012 20641 19014
rect 20697 19012 20721 19014
rect 20777 19012 20801 19014
rect 20857 19012 20863 19014
rect 20555 19003 20863 19012
rect 20916 18884 20944 19450
rect 22020 19310 22048 19790
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21192 18970 21220 19246
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 20824 18856 20944 18884
rect 20824 18766 20852 18856
rect 21284 18766 21312 18906
rect 22020 18766 22048 19110
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 20364 18426 20392 18634
rect 20916 18442 20944 18634
rect 20916 18426 21036 18442
rect 21468 18426 21496 18634
rect 22112 18426 22140 19314
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20352 18420 20404 18426
rect 20916 18420 21048 18426
rect 20916 18414 20996 18420
rect 20352 18362 20404 18368
rect 20996 18362 21048 18368
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 20272 18290 20300 18362
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20555 17980 20863 17989
rect 20555 17978 20561 17980
rect 20617 17978 20641 17980
rect 20697 17978 20721 17980
rect 20777 17978 20801 17980
rect 20857 17978 20863 17980
rect 20617 17926 20619 17978
rect 20799 17926 20801 17978
rect 20555 17924 20561 17926
rect 20617 17924 20641 17926
rect 20697 17924 20721 17926
rect 20777 17924 20801 17926
rect 20857 17924 20863 17926
rect 20555 17915 20863 17924
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19444 16658 19472 17138
rect 19536 17134 19564 17274
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19246 16552 19302 16561
rect 19246 16487 19302 16496
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 18880 15972 18932 15978
rect 18800 15932 18880 15960
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17420 13734 17448 14214
rect 17788 13802 17816 14962
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13870 18276 14214
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13326 17540 13670
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17788 13258 17816 13738
rect 18340 13410 18368 15302
rect 18524 15162 18552 15642
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18616 14958 18644 15302
rect 18708 14958 18736 15506
rect 18800 14958 18828 15932
rect 18880 15914 18932 15920
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19168 15366 19196 15506
rect 19260 15502 19288 15846
rect 19444 15552 19472 16458
rect 19536 15978 19564 17070
rect 19904 16998 19932 17818
rect 20916 17814 20944 18294
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19996 17270 20024 17478
rect 20272 17338 20300 17614
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 20732 17202 20760 17546
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 16250 19656 16390
rect 19720 16250 19748 16526
rect 19812 16522 19840 16934
rect 19996 16590 20024 17002
rect 20732 16998 20760 17138
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20555 16892 20863 16901
rect 20555 16890 20561 16892
rect 20617 16890 20641 16892
rect 20697 16890 20721 16892
rect 20777 16890 20801 16892
rect 20857 16890 20863 16892
rect 20617 16838 20619 16890
rect 20799 16838 20801 16890
rect 20555 16836 20561 16838
rect 20617 16836 20641 16838
rect 20697 16836 20721 16838
rect 20777 16836 20801 16838
rect 20857 16836 20863 16838
rect 20555 16827 20863 16836
rect 20916 16794 20944 17750
rect 21008 17241 21036 18362
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22020 18154 22048 18226
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 22112 18034 22140 18226
rect 22020 18006 22140 18034
rect 21086 17912 21142 17921
rect 21086 17847 21142 17856
rect 21100 17746 21128 17847
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 20994 17232 21050 17241
rect 20994 17167 21050 17176
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 21100 16726 21128 17546
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 21284 16658 21312 17138
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 21178 16552 21234 16561
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19628 15706 19656 16186
rect 19904 16046 19932 16390
rect 19996 16250 20024 16526
rect 20996 16516 21048 16522
rect 21178 16487 21180 16496
rect 20996 16458 21048 16464
rect 21232 16487 21234 16496
rect 21180 16458 21232 16464
rect 20076 16448 20128 16454
rect 21008 16425 21036 16458
rect 20076 16390 20128 16396
rect 20994 16416 21050 16425
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19996 16153 20024 16186
rect 19982 16144 20038 16153
rect 20088 16114 20116 16390
rect 20994 16351 21050 16360
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 19982 16079 20038 16088
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 20180 15570 20208 16186
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20555 15804 20863 15813
rect 20555 15802 20561 15804
rect 20617 15802 20641 15804
rect 20697 15802 20721 15804
rect 20777 15802 20801 15804
rect 20857 15802 20863 15804
rect 20617 15750 20619 15802
rect 20799 15750 20801 15802
rect 20555 15748 20561 15750
rect 20617 15748 20641 15750
rect 20697 15748 20721 15750
rect 20777 15748 20801 15750
rect 20857 15748 20863 15750
rect 20555 15739 20863 15748
rect 20916 15570 20944 16050
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20168 15564 20220 15570
rect 19444 15524 19564 15552
rect 19248 15496 19300 15502
rect 19536 15484 19564 15524
rect 20168 15506 20220 15512
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 19616 15496 19668 15502
rect 19536 15456 19616 15484
rect 19248 15438 19300 15444
rect 20444 15496 20496 15502
rect 19616 15438 19668 15444
rect 19982 15464 20038 15473
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 14958 19196 15302
rect 19260 15026 19288 15438
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 19156 14952 19208 14958
rect 19628 14940 19656 15438
rect 20444 15438 20496 15444
rect 19982 15399 20038 15408
rect 19708 14952 19760 14958
rect 19628 14912 19708 14940
rect 19156 14894 19208 14900
rect 19708 14894 19760 14900
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18432 13977 18460 14010
rect 18418 13968 18474 13977
rect 18418 13903 18474 13912
rect 18340 13394 18460 13410
rect 18340 13388 18472 13394
rect 18340 13382 18420 13388
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 18340 12986 18368 13382
rect 18420 13330 18472 13336
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16500 10062 16528 12378
rect 17132 12300 17184 12306
rect 17184 12260 17264 12288
rect 17132 12242 17184 12248
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 16634 11996 16942 12005
rect 16634 11994 16640 11996
rect 16696 11994 16720 11996
rect 16776 11994 16800 11996
rect 16856 11994 16880 11996
rect 16936 11994 16942 11996
rect 16696 11942 16698 11994
rect 16878 11942 16880 11994
rect 16634 11940 16640 11942
rect 16696 11940 16720 11942
rect 16776 11940 16800 11942
rect 16856 11940 16880 11942
rect 16936 11940 16942 11942
rect 16634 11931 16942 11940
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16868 11558 16896 11698
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 17052 11354 17080 12106
rect 17236 11762 17264 12260
rect 18248 12238 18276 12854
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18616 12170 18644 14894
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 11762 17816 12038
rect 17868 11824 17920 11830
rect 18800 11801 18828 14282
rect 18984 14278 19012 14894
rect 19996 14890 20024 15399
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18984 13530 19012 14214
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19524 13456 19576 13462
rect 19524 13398 19576 13404
rect 19444 12918 19472 13398
rect 19536 13190 19564 13398
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19536 12646 19564 13126
rect 19812 12782 19840 14350
rect 20180 13841 20208 14962
rect 20272 14822 20300 15302
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20364 14414 20392 15302
rect 20456 15026 20484 15438
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20824 15094 20852 15370
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20555 14716 20863 14725
rect 20555 14714 20561 14716
rect 20617 14714 20641 14716
rect 20697 14714 20721 14716
rect 20777 14714 20801 14716
rect 20857 14714 20863 14716
rect 20617 14662 20619 14714
rect 20799 14662 20801 14714
rect 20555 14660 20561 14662
rect 20617 14660 20641 14662
rect 20697 14660 20721 14662
rect 20777 14660 20801 14662
rect 20857 14660 20863 14662
rect 20555 14651 20863 14660
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20444 13864 20496 13870
rect 20166 13832 20222 13841
rect 20444 13806 20496 13812
rect 20166 13767 20222 13776
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 12986 20392 13262
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 20456 12714 20484 13806
rect 20555 13628 20863 13637
rect 20555 13626 20561 13628
rect 20617 13626 20641 13628
rect 20697 13626 20721 13628
rect 20777 13626 20801 13628
rect 20857 13626 20863 13628
rect 20617 13574 20619 13626
rect 20799 13574 20801 13626
rect 20555 13572 20561 13574
rect 20617 13572 20641 13574
rect 20697 13572 20721 13574
rect 20777 13572 20801 13574
rect 20857 13572 20863 13574
rect 20555 13563 20863 13572
rect 20916 12918 20944 15506
rect 21008 15502 21036 15846
rect 21100 15706 21128 15846
rect 21376 15706 21404 17138
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 21284 15201 21312 15506
rect 21270 15192 21326 15201
rect 21270 15127 21326 15136
rect 21468 15094 21496 17002
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21744 15638 21772 15982
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21640 15496 21692 15502
rect 21638 15464 21640 15473
rect 21692 15464 21694 15473
rect 21638 15399 21694 15408
rect 21732 15428 21784 15434
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21652 14958 21680 15399
rect 21732 15370 21784 15376
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21744 14618 21772 15370
rect 21836 14618 21864 15642
rect 21928 15337 21956 16594
rect 21914 15328 21970 15337
rect 21914 15263 21970 15272
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21744 13938 21772 14554
rect 21836 14278 21864 14554
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21928 13870 21956 15263
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21560 13326 21588 13466
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 21376 12850 21404 13126
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 20555 12540 20863 12549
rect 20555 12538 20561 12540
rect 20617 12538 20641 12540
rect 20697 12538 20721 12540
rect 20777 12538 20801 12540
rect 20857 12538 20863 12540
rect 20617 12486 20619 12538
rect 20799 12486 20801 12538
rect 20555 12484 20561 12486
rect 20617 12484 20641 12486
rect 20697 12484 20721 12486
rect 20777 12484 20801 12486
rect 20857 12484 20863 12486
rect 20555 12475 20863 12484
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 17868 11766 17920 11772
rect 18786 11792 18842 11801
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16946 11112 17002 11121
rect 17144 11082 17172 11494
rect 16946 11047 16948 11056
rect 17000 11047 17002 11056
rect 17132 11076 17184 11082
rect 16948 11018 17000 11024
rect 17132 11018 17184 11024
rect 16634 10908 16942 10917
rect 16634 10906 16640 10908
rect 16696 10906 16720 10908
rect 16776 10906 16800 10908
rect 16856 10906 16880 10908
rect 16936 10906 16942 10908
rect 16696 10854 16698 10906
rect 16878 10854 16880 10906
rect 16634 10852 16640 10854
rect 16696 10852 16720 10854
rect 16776 10852 16800 10854
rect 16856 10852 16880 10854
rect 16936 10852 16942 10854
rect 16634 10843 16942 10852
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16634 9820 16942 9829
rect 16634 9818 16640 9820
rect 16696 9818 16720 9820
rect 16776 9818 16800 9820
rect 16856 9818 16880 9820
rect 16936 9818 16942 9820
rect 16696 9766 16698 9818
rect 16878 9766 16880 9818
rect 16634 9764 16640 9766
rect 16696 9764 16720 9766
rect 16776 9764 16800 9766
rect 16856 9764 16880 9766
rect 16936 9764 16942 9766
rect 16634 9755 16942 9764
rect 17144 9654 17172 11018
rect 17236 10742 17264 11698
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17420 11354 17448 11630
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17788 11286 17816 11698
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17880 11150 17908 11766
rect 18786 11727 18788 11736
rect 18840 11727 18842 11736
rect 18972 11756 19024 11762
rect 18788 11698 18840 11704
rect 18972 11698 19024 11704
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17328 9926 17356 10542
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17328 9586 17356 9862
rect 17420 9654 17448 10950
rect 17972 10810 18000 11562
rect 18064 11218 18092 11630
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18984 10810 19012 11698
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11286 19104 11494
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19168 10742 19196 12038
rect 19444 11354 19472 12174
rect 20555 11452 20863 11461
rect 20555 11450 20561 11452
rect 20617 11450 20641 11452
rect 20697 11450 20721 11452
rect 20777 11450 20801 11452
rect 20857 11450 20863 11452
rect 20617 11398 20619 11450
rect 20799 11398 20801 11450
rect 20555 11396 20561 11398
rect 20617 11396 20641 11398
rect 20697 11396 20721 11398
rect 20777 11396 20801 11398
rect 20857 11396 20863 11398
rect 20555 11387 20863 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9926 17540 10066
rect 18248 9994 18276 10542
rect 18340 10062 18368 10610
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18432 10010 18460 10202
rect 18524 10198 18552 10610
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 18616 10010 18644 10202
rect 18800 10198 18828 10474
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8498 16252 8774
rect 16634 8732 16942 8741
rect 16634 8730 16640 8732
rect 16696 8730 16720 8732
rect 16776 8730 16800 8732
rect 16856 8730 16880 8732
rect 16936 8730 16942 8732
rect 16696 8678 16698 8730
rect 16878 8678 16880 8730
rect 16634 8676 16640 8678
rect 16696 8676 16720 8678
rect 16776 8676 16800 8678
rect 16856 8676 16880 8678
rect 16936 8676 16942 8678
rect 16634 8667 16942 8676
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 17052 8090 17080 8910
rect 17144 8906 17172 9318
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 16408 7546 16436 7754
rect 16634 7644 16942 7653
rect 16634 7642 16640 7644
rect 16696 7642 16720 7644
rect 16776 7642 16800 7644
rect 16856 7642 16880 7644
rect 16936 7642 16942 7644
rect 16696 7590 16698 7642
rect 16878 7590 16880 7642
rect 16634 7588 16640 7590
rect 16696 7588 16720 7590
rect 16776 7588 16800 7590
rect 16856 7588 16880 7590
rect 16936 7588 16942 7590
rect 16634 7579 16942 7588
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 17052 6882 17080 7890
rect 17144 7886 17172 8842
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8294 17264 8774
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17236 7732 17264 8230
rect 17328 7886 17356 9386
rect 17512 8650 17540 9862
rect 18248 9586 18276 9930
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 9178 18276 9522
rect 18340 9450 18368 9998
rect 18432 9982 18644 10010
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 17420 8622 17540 8650
rect 17420 8022 17448 8622
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17512 8090 17540 8434
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17236 7704 17356 7732
rect 17328 7342 17356 7704
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16960 6854 17080 6882
rect 14844 6322 14872 6802
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6322 15884 6734
rect 16132 6322 16160 6802
rect 16960 6798 16988 6854
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16634 6556 16942 6565
rect 16634 6554 16640 6556
rect 16696 6554 16720 6556
rect 16776 6554 16800 6556
rect 16856 6554 16880 6556
rect 16936 6554 16942 6556
rect 16696 6502 16698 6554
rect 16878 6502 16880 6554
rect 16634 6500 16640 6502
rect 16696 6500 16720 6502
rect 16776 6500 16800 6502
rect 16856 6500 16880 6502
rect 16936 6500 16942 6502
rect 16634 6491 16942 6500
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 14844 5710 14872 6258
rect 16500 6118 16528 6258
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16224 5778 16252 6054
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 8792 5468 9100 5477
rect 8792 5466 8798 5468
rect 8854 5466 8878 5468
rect 8934 5466 8958 5468
rect 9014 5466 9038 5468
rect 9094 5466 9100 5468
rect 8854 5414 8856 5466
rect 9036 5414 9038 5466
rect 8792 5412 8798 5414
rect 8854 5412 8878 5414
rect 8934 5412 8958 5414
rect 9014 5412 9038 5414
rect 9094 5412 9100 5414
rect 8792 5403 9100 5412
rect 16634 5468 16942 5477
rect 16634 5466 16640 5468
rect 16696 5466 16720 5468
rect 16776 5466 16800 5468
rect 16856 5466 16880 5468
rect 16936 5466 16942 5468
rect 16696 5414 16698 5466
rect 16878 5414 16880 5466
rect 16634 5412 16640 5414
rect 16696 5412 16720 5414
rect 16776 5412 16800 5414
rect 16856 5412 16880 5414
rect 16936 5412 16942 5414
rect 16634 5403 16942 5412
rect 17052 5370 17080 6734
rect 17144 6458 17172 7142
rect 17236 7002 17264 7278
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17604 6866 17632 9046
rect 18524 8906 18552 9046
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18524 8566 18552 8842
rect 18616 8634 18644 9982
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9586 19288 9862
rect 19352 9654 19380 10542
rect 19536 10266 19564 10542
rect 19628 10266 19656 10950
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19536 9586 19564 10202
rect 19812 9926 19840 10610
rect 20180 10470 20208 11018
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19812 9722 19840 9862
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 9178 19380 9454
rect 19444 9178 19472 9522
rect 19628 9382 19656 9590
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17696 7546 17724 7754
rect 17880 7546 17908 7822
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18616 7410 18644 8570
rect 18708 8498 18736 8774
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 7002 18000 7210
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5914 17172 6190
rect 17236 6186 17264 6734
rect 17328 6322 17356 6802
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17144 5642 17172 5850
rect 17236 5710 17264 6122
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17144 5302 17172 5578
rect 17328 5574 17356 6258
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17512 5778 17540 6190
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17512 5234 17540 5714
rect 17604 5710 17632 6802
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6118 18184 6598
rect 18616 6322 18644 7346
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5846 18184 6054
rect 18616 5914 18644 6258
rect 19352 6186 19380 9114
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19444 7954 19472 8774
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19628 7886 19656 8774
rect 19904 8090 19932 8842
rect 20272 8634 20300 11086
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10062 20392 10406
rect 20555 10364 20863 10373
rect 20555 10362 20561 10364
rect 20617 10362 20641 10364
rect 20697 10362 20721 10364
rect 20777 10362 20801 10364
rect 20857 10362 20863 10364
rect 20617 10310 20619 10362
rect 20799 10310 20801 10362
rect 20555 10308 20561 10310
rect 20617 10308 20641 10310
rect 20697 10308 20721 10310
rect 20777 10308 20801 10310
rect 20857 10308 20863 10310
rect 20555 10299 20863 10308
rect 20916 10130 20944 12718
rect 21560 12442 21588 13262
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21928 10538 21956 13806
rect 22020 13433 22048 18006
rect 22204 17320 22232 19382
rect 22296 19310 22324 19790
rect 22284 19304 22336 19310
rect 22282 19272 22284 19281
rect 22336 19272 22338 19281
rect 22282 19207 22338 19216
rect 22388 18902 22416 19858
rect 23032 19854 23060 20266
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22560 18284 22612 18290
rect 22664 18272 22692 19110
rect 22756 18426 22784 19246
rect 23216 18766 23244 19314
rect 23584 18902 23612 20402
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24476 19612 24784 19621
rect 24476 19610 24482 19612
rect 24538 19610 24562 19612
rect 24618 19610 24642 19612
rect 24698 19610 24722 19612
rect 24778 19610 24784 19612
rect 24538 19558 24540 19610
rect 24720 19558 24722 19610
rect 24476 19556 24482 19558
rect 24538 19556 24562 19558
rect 24618 19556 24642 19558
rect 24698 19556 24722 19558
rect 24778 19556 24784 19558
rect 24476 19547 24784 19556
rect 24872 19242 24900 19858
rect 24964 19854 24992 20198
rect 25976 19938 26004 20334
rect 25884 19910 26004 19938
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25884 19446 25912 19910
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25872 19440 25924 19446
rect 25872 19382 25924 19388
rect 25884 19242 25912 19382
rect 25976 19310 26004 19654
rect 26252 19378 26280 20402
rect 27816 20058 27844 20402
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26712 19514 26740 19790
rect 26804 19514 26832 19858
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 27896 19712 27948 19718
rect 27896 19654 27948 19660
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 26252 18902 26280 19314
rect 26424 19304 26476 19310
rect 26424 19246 26476 19252
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 26240 18896 26292 18902
rect 26240 18838 26292 18844
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22744 18284 22796 18290
rect 22612 18244 22744 18272
rect 22560 18226 22612 18232
rect 22744 18226 22796 18232
rect 23216 17882 23244 18702
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23400 18426 23428 18566
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 24412 18290 24440 18702
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24476 18524 24784 18533
rect 24476 18522 24482 18524
rect 24538 18522 24562 18524
rect 24618 18522 24642 18524
rect 24698 18522 24722 18524
rect 24778 18522 24784 18524
rect 24538 18470 24540 18522
rect 24720 18470 24722 18522
rect 24476 18468 24482 18470
rect 24538 18468 24562 18470
rect 24618 18468 24642 18470
rect 24698 18468 24722 18470
rect 24778 18468 24784 18470
rect 24476 18459 24784 18468
rect 24872 18290 24900 18634
rect 25148 18290 25176 18702
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 22204 17292 22324 17320
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 16590 22140 16934
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22204 15162 22232 17138
rect 22296 16454 22324 17292
rect 23124 17134 23152 17682
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23308 17542 23336 17614
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23400 17270 23428 18022
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23492 17338 23520 17546
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23124 16794 23152 17070
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22190 14920 22246 14929
rect 22190 14855 22246 14864
rect 22204 14482 22232 14855
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22192 13932 22244 13938
rect 22296 13920 22324 15438
rect 22756 15434 22784 15846
rect 22940 15570 22968 15846
rect 23216 15706 23244 16118
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22244 13892 22324 13920
rect 22192 13874 22244 13880
rect 22006 13424 22062 13433
rect 22006 13359 22062 13368
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22112 12170 22140 12718
rect 22204 12646 22232 13874
rect 22388 13870 22416 14962
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22480 14414 22508 14758
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22204 11762 22232 12582
rect 22296 12306 22324 12650
rect 22388 12434 22416 13670
rect 22572 13546 22600 14418
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22664 13734 22692 14350
rect 22940 13870 22968 15506
rect 23216 15026 23244 15506
rect 23480 15496 23532 15502
rect 23478 15464 23480 15473
rect 23532 15464 23534 15473
rect 23478 15399 23534 15408
rect 23584 15094 23612 17750
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23676 16561 23704 17546
rect 23662 16552 23718 16561
rect 23662 16487 23718 16496
rect 23768 16153 23796 17818
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23754 16144 23810 16153
rect 23754 16079 23810 16088
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23676 15570 23704 15914
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23676 15337 23704 15506
rect 23768 15502 23796 16079
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23662 15328 23718 15337
rect 23662 15263 23718 15272
rect 23662 15192 23718 15201
rect 23662 15127 23718 15136
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23308 14618 23336 14962
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23124 13938 23152 14418
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22572 13518 22692 13546
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22388 12406 22508 12434
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22020 10674 22048 10746
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20916 9466 20944 10066
rect 21928 9654 21956 10474
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 20456 8906 20484 9454
rect 20916 9450 21128 9466
rect 20916 9444 21140 9450
rect 20916 9438 21088 9444
rect 20555 9276 20863 9285
rect 20555 9274 20561 9276
rect 20617 9274 20641 9276
rect 20697 9274 20721 9276
rect 20777 9274 20801 9276
rect 20857 9274 20863 9276
rect 20617 9222 20619 9274
rect 20799 9222 20801 9274
rect 20555 9220 20561 9222
rect 20617 9220 20641 9222
rect 20697 9220 20721 9222
rect 20777 9220 20801 9222
rect 20857 9220 20863 9222
rect 20555 9211 20863 9220
rect 20718 9072 20774 9081
rect 20718 9007 20774 9016
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19536 7546 19564 7822
rect 20272 7750 20300 8570
rect 20732 8498 20760 9007
rect 20916 8974 20944 9438
rect 21088 9386 21140 9392
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 21928 8974 21956 9386
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21364 8900 21416 8906
rect 21364 8842 21416 8848
rect 21376 8566 21404 8842
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21928 8498 21956 8910
rect 22020 8838 22048 10610
rect 22204 9722 22232 10610
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22388 8634 22416 11290
rect 22480 10606 22508 12406
rect 22572 12306 22600 13330
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22572 11626 22600 12242
rect 22664 12102 22692 13518
rect 23308 13258 23336 14554
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22756 12850 22784 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22756 12238 22784 12786
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 12442 22876 12582
rect 23216 12442 23244 12718
rect 23308 12646 23336 12922
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23308 12374 23336 12582
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22480 8974 22508 10406
rect 22572 9654 22600 10610
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 20555 8188 20863 8197
rect 20555 8186 20561 8188
rect 20617 8186 20641 8188
rect 20697 8186 20721 8188
rect 20777 8186 20801 8188
rect 20857 8186 20863 8188
rect 20617 8134 20619 8186
rect 20799 8134 20801 8186
rect 20555 8132 20561 8134
rect 20617 8132 20641 8134
rect 20697 8132 20721 8134
rect 20777 8132 20801 8134
rect 20857 8132 20863 8134
rect 20555 8123 20863 8132
rect 21192 8090 21220 8434
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 22388 7954 22416 8570
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 20272 7274 20300 7686
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 20444 7336 20496 7342
rect 20364 7284 20444 7290
rect 20364 7278 20496 7284
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20364 7262 20484 7278
rect 20364 6798 20392 7262
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 20456 7002 20484 7142
rect 20555 7100 20863 7109
rect 20555 7098 20561 7100
rect 20617 7098 20641 7100
rect 20697 7098 20721 7100
rect 20777 7098 20801 7100
rect 20857 7098 20863 7100
rect 20617 7046 20619 7098
rect 20799 7046 20801 7098
rect 20555 7044 20561 7046
rect 20617 7044 20641 7046
rect 20697 7044 20721 7046
rect 20777 7044 20801 7046
rect 20857 7044 20863 7046
rect 20555 7035 20863 7044
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20812 6928 20864 6934
rect 20812 6870 20864 6876
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 19628 6390 19656 6734
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20088 6458 20116 6598
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19616 6384 19668 6390
rect 19616 6326 19668 6332
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 19628 5234 19656 6326
rect 20824 6322 20852 6870
rect 20904 6792 20956 6798
rect 21088 6792 21140 6798
rect 20956 6752 21036 6780
rect 20904 6734 20956 6740
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20272 5778 20300 6122
rect 20456 5846 20484 6122
rect 20555 6012 20863 6021
rect 20555 6010 20561 6012
rect 20617 6010 20641 6012
rect 20697 6010 20721 6012
rect 20777 6010 20801 6012
rect 20857 6010 20863 6012
rect 20617 5958 20619 6010
rect 20799 5958 20801 6010
rect 20555 5956 20561 5958
rect 20617 5956 20641 5958
rect 20697 5956 20721 5958
rect 20777 5956 20801 5958
rect 20857 5956 20863 5958
rect 20555 5947 20863 5956
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 20272 5030 20300 5714
rect 20916 5370 20944 6122
rect 21008 5914 21036 6752
rect 21088 6734 21140 6740
rect 21100 6662 21128 6734
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6322 21128 6598
rect 21192 6322 21220 7142
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21100 5914 21128 6258
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 21100 5234 21128 5714
rect 21376 5234 21404 6870
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21468 6254 21496 6734
rect 21560 6458 21588 6734
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21560 5846 21588 6394
rect 21652 5914 21680 7482
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21744 6934 21772 7142
rect 22388 6934 22416 7754
rect 22572 7410 22600 7890
rect 22664 7478 22692 12038
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22756 11150 22784 11494
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23124 10266 23152 11086
rect 23400 10742 23428 14010
rect 23676 13546 23704 15127
rect 23492 13518 23704 13546
rect 23492 10810 23520 13518
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23676 12170 23704 12922
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23676 11218 23704 11766
rect 23768 11286 23796 15438
rect 23860 14770 23888 16526
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23952 15570 23980 16390
rect 24044 16250 24072 18226
rect 24872 17678 24900 18226
rect 25148 17882 25176 18226
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 25148 17785 25176 17818
rect 25134 17776 25190 17785
rect 25134 17711 25190 17720
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24320 16794 24348 17478
rect 24476 17436 24784 17445
rect 24476 17434 24482 17436
rect 24538 17434 24562 17436
rect 24618 17434 24642 17436
rect 24698 17434 24722 17436
rect 24778 17434 24784 17436
rect 24538 17382 24540 17434
rect 24720 17382 24722 17434
rect 24476 17380 24482 17382
rect 24538 17380 24562 17382
rect 24618 17380 24642 17382
rect 24698 17380 24722 17382
rect 24778 17380 24784 17382
rect 24476 17371 24784 17380
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24136 16182 24164 16526
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 24320 15978 24348 16730
rect 24780 16590 24808 17138
rect 24964 17066 24992 17546
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 25240 16794 25268 18022
rect 25976 17921 26004 18566
rect 25962 17912 26018 17921
rect 25962 17847 26018 17856
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25516 16998 25544 17138
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24214 15192 24270 15201
rect 24214 15127 24216 15136
rect 24268 15127 24270 15136
rect 24216 15098 24268 15104
rect 23940 14816 23992 14822
rect 23860 14764 23940 14770
rect 23860 14758 23992 14764
rect 23860 14742 23980 14758
rect 23860 14278 23888 14742
rect 24320 14618 24348 15302
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24228 13938 24256 14214
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24320 13870 24348 14554
rect 24412 14414 24440 16390
rect 24476 16348 24784 16357
rect 24476 16346 24482 16348
rect 24538 16346 24562 16348
rect 24618 16346 24642 16348
rect 24698 16346 24722 16348
rect 24778 16346 24784 16348
rect 24538 16294 24540 16346
rect 24720 16294 24722 16346
rect 24476 16292 24482 16294
rect 24538 16292 24562 16294
rect 24618 16292 24642 16294
rect 24698 16292 24722 16294
rect 24778 16292 24784 16294
rect 24476 16283 24784 16292
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24476 15260 24784 15269
rect 24476 15258 24482 15260
rect 24538 15258 24562 15260
rect 24618 15258 24642 15260
rect 24698 15258 24722 15260
rect 24778 15258 24784 15260
rect 24538 15206 24540 15258
rect 24720 15206 24722 15258
rect 24476 15204 24482 15206
rect 24538 15204 24562 15206
rect 24618 15204 24642 15206
rect 24698 15204 24722 15206
rect 24778 15204 24784 15206
rect 24476 15195 24784 15204
rect 24872 15026 24900 15370
rect 24964 15162 24992 15846
rect 25056 15706 25084 16050
rect 25148 15978 25176 16594
rect 25240 16522 25268 16730
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 25136 15972 25188 15978
rect 25136 15914 25188 15920
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 25240 15502 25268 16458
rect 25608 16250 25636 17138
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25332 15502 25360 15642
rect 25424 15502 25452 16050
rect 25700 15502 25728 17002
rect 25792 15638 25820 17478
rect 25872 16040 25924 16046
rect 25870 16008 25872 16017
rect 25924 16008 25926 16017
rect 25870 15943 25926 15952
rect 25780 15632 25832 15638
rect 25780 15574 25832 15580
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25320 15496 25372 15502
rect 25412 15496 25464 15502
rect 25320 15438 25372 15444
rect 25410 15464 25412 15473
rect 25688 15496 25740 15502
rect 25464 15464 25466 15473
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24964 14414 24992 15098
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25148 14618 25176 15030
rect 25240 14618 25268 15438
rect 25466 15422 25636 15450
rect 25688 15438 25740 15444
rect 25410 15399 25466 15408
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25136 14612 25188 14618
rect 25056 14572 25136 14600
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24412 13938 24440 14350
rect 24964 14278 24992 14350
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24476 14172 24784 14181
rect 24476 14170 24482 14172
rect 24538 14170 24562 14172
rect 24618 14170 24642 14172
rect 24698 14170 24722 14172
rect 24778 14170 24784 14172
rect 24538 14118 24540 14170
rect 24720 14118 24722 14170
rect 24476 14116 24482 14118
rect 24538 14116 24562 14118
rect 24618 14116 24642 14118
rect 24698 14116 24722 14118
rect 24778 14116 24784 14118
rect 24476 14107 24784 14116
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 25056 13870 25084 14572
rect 25136 14554 25188 14560
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 24308 13864 24360 13870
rect 24214 13832 24270 13841
rect 24308 13806 24360 13812
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 24214 13767 24270 13776
rect 24228 13734 24256 13767
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24228 13326 24256 13670
rect 24308 13388 24360 13394
rect 24308 13330 24360 13336
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23860 12850 23888 13126
rect 24320 12850 24348 13330
rect 24674 13288 24730 13297
rect 24674 13223 24676 13232
rect 24728 13223 24730 13232
rect 24676 13194 24728 13200
rect 24476 13084 24784 13093
rect 24476 13082 24482 13084
rect 24538 13082 24562 13084
rect 24618 13082 24642 13084
rect 24698 13082 24722 13084
rect 24778 13082 24784 13084
rect 24538 13030 24540 13082
rect 24720 13030 24722 13082
rect 24476 13028 24482 13030
rect 24538 13028 24562 13030
rect 24618 13028 24642 13030
rect 24698 13028 24722 13030
rect 24778 13028 24784 13030
rect 24476 13019 24784 13028
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 23860 11694 23888 12786
rect 24688 12374 24716 12922
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 24964 12238 24992 12922
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24476 11996 24784 12005
rect 24476 11994 24482 11996
rect 24538 11994 24562 11996
rect 24618 11994 24642 11996
rect 24698 11994 24722 11996
rect 24778 11994 24784 11996
rect 24538 11942 24540 11994
rect 24720 11942 24722 11994
rect 24476 11940 24482 11942
rect 24538 11940 24562 11942
rect 24618 11940 24642 11942
rect 24698 11940 24722 11942
rect 24778 11940 24784 11942
rect 24476 11931 24784 11940
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23952 11354 23980 11698
rect 25148 11354 25176 14350
rect 25332 14278 25360 14758
rect 25412 14340 25464 14346
rect 25412 14282 25464 14288
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25240 12986 25268 13874
rect 25332 13734 25360 14214
rect 25424 13938 25452 14282
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25332 13326 25360 13670
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 25516 12306 25544 12854
rect 25608 12782 25636 15422
rect 25976 15026 26004 17847
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 26068 17338 26096 17614
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 26068 16658 26096 17274
rect 26160 16998 26188 18702
rect 26344 18290 26372 19110
rect 26436 18426 26464 19246
rect 26528 18970 26556 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 27356 18766 27384 19110
rect 27448 18970 27476 19382
rect 27908 19378 27936 19654
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 28092 18970 28120 19790
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 27448 18290 27476 18906
rect 28276 18766 28304 21383
rect 28397 20156 28705 20165
rect 28397 20154 28403 20156
rect 28459 20154 28483 20156
rect 28539 20154 28563 20156
rect 28619 20154 28643 20156
rect 28699 20154 28705 20156
rect 28459 20102 28461 20154
rect 28641 20102 28643 20154
rect 28397 20100 28403 20102
rect 28459 20100 28483 20102
rect 28539 20100 28563 20102
rect 28619 20100 28643 20102
rect 28699 20100 28705 20102
rect 28397 20091 28705 20100
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28368 19514 28396 19790
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28397 19068 28705 19077
rect 28397 19066 28403 19068
rect 28459 19066 28483 19068
rect 28539 19066 28563 19068
rect 28619 19066 28643 19068
rect 28699 19066 28705 19068
rect 28459 19014 28461 19066
rect 28641 19014 28643 19066
rect 28397 19012 28403 19014
rect 28459 19012 28483 19014
rect 28539 19012 28563 19014
rect 28619 19012 28643 19014
rect 28699 19012 28705 19014
rect 28397 19003 28705 19012
rect 28736 18766 28764 21383
rect 29184 20256 29236 20262
rect 29184 20198 29236 20204
rect 29196 19514 29224 20198
rect 29472 19990 29500 21383
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29460 19984 29512 19990
rect 29460 19926 29512 19932
rect 29748 19854 29776 20334
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 28816 19440 28868 19446
rect 28816 19382 28868 19388
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26330 17640 26386 17649
rect 26330 17575 26386 17584
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26252 17338 26280 17478
rect 26344 17338 26372 17575
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26068 15502 26096 16458
rect 26252 16454 26280 17138
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 25780 15020 25832 15026
rect 25780 14962 25832 14968
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25700 12850 25728 14758
rect 25792 14482 25820 14962
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25884 14414 25912 14894
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25962 14376 26018 14385
rect 25884 13870 25912 14350
rect 25962 14311 25964 14320
rect 26016 14311 26018 14320
rect 25964 14282 26016 14288
rect 26068 14074 26096 15438
rect 26252 15162 26280 16390
rect 26344 16114 26372 17274
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26436 16658 26464 17138
rect 26528 16794 26556 17682
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26620 17338 26648 17546
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 27264 17134 27292 18022
rect 27448 17542 27476 18226
rect 28397 17980 28705 17989
rect 28397 17978 28403 17980
rect 28459 17978 28483 17980
rect 28539 17978 28563 17980
rect 28619 17978 28643 17980
rect 28699 17978 28705 17980
rect 28459 17926 28461 17978
rect 28641 17926 28643 17978
rect 28397 17924 28403 17926
rect 28459 17924 28483 17926
rect 28539 17924 28563 17926
rect 28619 17924 28643 17926
rect 28699 17924 28705 17926
rect 28397 17915 28705 17924
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 27436 17536 27488 17542
rect 27436 17478 27488 17484
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 26516 16788 26568 16794
rect 26516 16730 26568 16736
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26436 16017 26464 16594
rect 27632 16182 27660 16934
rect 28276 16726 28304 17138
rect 28397 16892 28705 16901
rect 28397 16890 28403 16892
rect 28459 16890 28483 16892
rect 28539 16890 28563 16892
rect 28619 16890 28643 16892
rect 28699 16890 28705 16892
rect 28459 16838 28461 16890
rect 28641 16838 28643 16890
rect 28397 16836 28403 16838
rect 28459 16836 28483 16838
rect 28539 16836 28563 16838
rect 28619 16836 28643 16838
rect 28699 16836 28705 16838
rect 28397 16827 28705 16836
rect 28264 16720 28316 16726
rect 28264 16662 28316 16668
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 26608 16176 26660 16182
rect 26608 16118 26660 16124
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 26422 16008 26478 16017
rect 26422 15943 26478 15952
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 26252 14521 26280 14554
rect 26344 14550 26372 14962
rect 26332 14544 26384 14550
rect 26238 14512 26294 14521
rect 26332 14486 26384 14492
rect 26238 14447 26294 14456
rect 26240 14408 26292 14414
rect 26160 14356 26240 14362
rect 26160 14350 26292 14356
rect 26160 14334 26280 14350
rect 26160 14278 26188 14334
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25608 12322 25636 12718
rect 25504 12300 25556 12306
rect 25608 12294 25728 12322
rect 25504 12242 25556 12248
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23952 11150 23980 11290
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 23216 9994 23244 10134
rect 23204 9988 23256 9994
rect 23204 9930 23256 9936
rect 23308 7818 23336 10610
rect 23400 10130 23428 10678
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23492 9042 23520 10746
rect 23676 10266 23704 11018
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24476 10908 24784 10917
rect 24476 10906 24482 10908
rect 24538 10906 24562 10908
rect 24618 10906 24642 10908
rect 24698 10906 24722 10908
rect 24778 10906 24784 10908
rect 24538 10854 24540 10906
rect 24720 10854 24722 10906
rect 24476 10852 24482 10854
rect 24538 10852 24562 10854
rect 24618 10852 24642 10854
rect 24698 10852 24722 10854
rect 24778 10852 24784 10854
rect 24476 10843 24784 10852
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23676 9654 23704 9930
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23676 8838 23704 9590
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23492 8022 23520 8434
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23584 8090 23612 8230
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 21744 6798 21772 6870
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 21744 5574 21772 6190
rect 21836 5710 21864 6598
rect 22480 6322 22508 7210
rect 22572 6866 22600 7346
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 23032 6798 23060 7278
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22480 5914 22508 6258
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 23032 5710 23060 6734
rect 23308 6662 23336 7754
rect 23676 7274 23704 8774
rect 24320 8634 24348 9522
rect 24412 8634 24440 10406
rect 24964 10062 24992 10950
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24476 9820 24784 9829
rect 24476 9818 24482 9820
rect 24538 9818 24562 9820
rect 24618 9818 24642 9820
rect 24698 9818 24722 9820
rect 24778 9818 24784 9820
rect 24538 9766 24540 9818
rect 24720 9766 24722 9818
rect 24476 9764 24482 9766
rect 24538 9764 24562 9766
rect 24618 9764 24642 9766
rect 24698 9764 24722 9766
rect 24778 9764 24784 9766
rect 24476 9755 24784 9764
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24780 8974 24808 9318
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24476 8732 24784 8741
rect 24476 8730 24482 8732
rect 24538 8730 24562 8732
rect 24618 8730 24642 8732
rect 24698 8730 24722 8732
rect 24778 8730 24784 8732
rect 24538 8678 24540 8730
rect 24720 8678 24722 8730
rect 24476 8676 24482 8678
rect 24538 8676 24562 8678
rect 24618 8676 24642 8678
rect 24698 8676 24722 8678
rect 24778 8676 24784 8678
rect 24476 8667 24784 8676
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24872 8498 24900 9862
rect 24964 9518 24992 9998
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25056 9722 25084 9862
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 25332 9654 25360 12038
rect 25608 10810 25636 12174
rect 25700 12170 25728 12294
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25700 11830 25728 12106
rect 25792 11898 25820 12174
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25688 11824 25740 11830
rect 25688 11766 25740 11772
rect 25884 11354 25912 13670
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 25976 13258 26004 13466
rect 26148 13456 26200 13462
rect 26068 13416 26148 13444
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 26068 12850 26096 13416
rect 26148 13398 26200 13404
rect 26252 13394 26280 14214
rect 26528 13938 26556 14962
rect 26620 14822 26648 16118
rect 28184 16114 28212 16458
rect 28644 16250 28672 16458
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28184 15910 28212 16050
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28397 15804 28705 15813
rect 28397 15802 28403 15804
rect 28459 15802 28483 15804
rect 28539 15802 28563 15804
rect 28619 15802 28643 15804
rect 28699 15802 28705 15804
rect 28459 15750 28461 15802
rect 28641 15750 28643 15802
rect 28397 15748 28403 15750
rect 28459 15748 28483 15750
rect 28539 15748 28563 15750
rect 28619 15748 28643 15750
rect 28699 15748 28705 15750
rect 28397 15739 28705 15748
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 26792 15632 26844 15638
rect 26792 15574 26844 15580
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26344 13394 26372 13466
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26528 13326 26556 13874
rect 26620 13802 26648 14418
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26608 13796 26660 13802
rect 26608 13738 26660 13744
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26160 12986 26188 13194
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25976 12306 26004 12718
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 25976 11830 26004 12242
rect 26068 12238 26096 12786
rect 26252 12442 26280 13194
rect 26240 12436 26292 12442
rect 26240 12378 26292 12384
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25884 11150 25912 11290
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 25424 9081 25452 9998
rect 25410 9072 25466 9081
rect 25410 9007 25466 9016
rect 25792 8838 25820 11086
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 26068 10062 26096 10950
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 26608 10736 26660 10742
rect 26712 10724 26740 13806
rect 26804 13326 26832 15574
rect 27448 15366 27476 15642
rect 28552 15366 28580 15642
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27712 15360 27764 15366
rect 27712 15302 27764 15308
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 27448 15094 27476 15302
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27448 14414 27476 15030
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27540 13410 27568 14758
rect 27724 14482 27752 15302
rect 28736 15162 28764 17614
rect 28828 17134 28856 19382
rect 30300 18698 30328 19790
rect 30484 18970 30512 20402
rect 31668 20256 31720 20262
rect 31668 20198 31720 20204
rect 30932 19848 30984 19854
rect 30932 19790 30984 19796
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30944 18698 30972 19790
rect 31576 19712 31628 19718
rect 31576 19654 31628 19660
rect 31484 19508 31536 19514
rect 31484 19450 31536 19456
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 30932 18692 30984 18698
rect 30932 18634 30984 18640
rect 29184 18624 29236 18630
rect 29184 18566 29236 18572
rect 29196 18290 29224 18566
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 29104 17134 29132 18158
rect 30300 17678 30328 18634
rect 30380 18080 30432 18086
rect 30380 18022 30432 18028
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 29736 17604 29788 17610
rect 29736 17546 29788 17552
rect 28816 17128 28868 17134
rect 28816 17070 28868 17076
rect 29092 17128 29144 17134
rect 29092 17070 29144 17076
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28080 15088 28132 15094
rect 28080 15030 28132 15036
rect 28264 15088 28316 15094
rect 28264 15030 28316 15036
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27724 13938 27752 14418
rect 28092 14278 28120 15030
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28184 14618 28212 14758
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27816 13530 27844 13874
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27540 13382 27844 13410
rect 27816 13326 27844 13382
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 26660 10696 26740 10724
rect 26608 10678 26660 10684
rect 26332 10532 26384 10538
rect 26332 10474 26384 10480
rect 26344 10062 26372 10474
rect 26528 10062 26556 10678
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26332 10056 26384 10062
rect 26332 9998 26384 10004
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25976 8974 26004 9862
rect 26068 9722 26096 9998
rect 26620 9994 26648 10678
rect 26804 10198 26832 13262
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27448 12986 27476 13126
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 26792 10192 26844 10198
rect 26792 10134 26844 10140
rect 26608 9988 26660 9994
rect 26608 9930 26660 9936
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 26528 9710 26740 9738
rect 26148 9648 26200 9654
rect 26148 9590 26200 9596
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 26160 9450 26188 9590
rect 26148 9444 26200 9450
rect 26148 9386 26200 9392
rect 26160 9110 26188 9386
rect 26252 9382 26280 9590
rect 26528 9382 26556 9710
rect 26712 9654 26740 9710
rect 27264 9654 27292 12786
rect 27632 12714 27660 13262
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27724 12850 27752 13126
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27620 12708 27672 12714
rect 27620 12650 27672 12656
rect 27724 12442 27752 12786
rect 27908 12782 27936 13126
rect 27896 12776 27948 12782
rect 27896 12718 27948 12724
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 27908 11762 27936 12718
rect 27988 12708 28040 12714
rect 27988 12650 28040 12656
rect 28000 11762 28028 12650
rect 28092 12434 28120 14214
rect 28276 13530 28304 15030
rect 28397 14716 28705 14725
rect 28397 14714 28403 14716
rect 28459 14714 28483 14716
rect 28539 14714 28563 14716
rect 28619 14714 28643 14716
rect 28699 14714 28705 14716
rect 28459 14662 28461 14714
rect 28641 14662 28643 14714
rect 28397 14660 28403 14662
rect 28459 14660 28483 14662
rect 28539 14660 28563 14662
rect 28619 14660 28643 14662
rect 28699 14660 28705 14662
rect 28397 14651 28705 14660
rect 28722 14512 28778 14521
rect 28828 14482 28856 17070
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28920 16114 28948 16934
rect 29104 16794 29132 17070
rect 29092 16788 29144 16794
rect 29092 16730 29144 16736
rect 29748 16250 29776 17546
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 29840 16590 29868 17478
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29736 16244 29788 16250
rect 29736 16186 29788 16192
rect 28908 16108 28960 16114
rect 28908 16050 28960 16056
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29288 15706 29316 15982
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 28908 14952 28960 14958
rect 28908 14894 28960 14900
rect 28722 14447 28778 14456
rect 28816 14476 28868 14482
rect 28736 14278 28764 14447
rect 28816 14418 28868 14424
rect 28920 14414 28948 14894
rect 28908 14408 28960 14414
rect 28814 14376 28870 14385
rect 28908 14350 28960 14356
rect 28814 14311 28816 14320
rect 28868 14311 28870 14320
rect 28816 14282 28868 14288
rect 28724 14272 28776 14278
rect 28724 14214 28776 14220
rect 28397 13628 28705 13637
rect 28397 13626 28403 13628
rect 28459 13626 28483 13628
rect 28539 13626 28563 13628
rect 28619 13626 28643 13628
rect 28699 13626 28705 13628
rect 28459 13574 28461 13626
rect 28641 13574 28643 13626
rect 28397 13572 28403 13574
rect 28459 13572 28483 13574
rect 28539 13572 28563 13574
rect 28619 13572 28643 13574
rect 28699 13572 28705 13574
rect 28397 13563 28705 13572
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 28736 13326 28764 14214
rect 28920 14006 28948 14350
rect 28908 14000 28960 14006
rect 28908 13942 28960 13948
rect 29012 13462 29040 15438
rect 29736 15156 29788 15162
rect 29736 15098 29788 15104
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29380 13938 29408 14962
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29368 13932 29420 13938
rect 29368 13874 29420 13880
rect 29092 13728 29144 13734
rect 29092 13670 29144 13676
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 29000 13320 29052 13326
rect 29104 13274 29132 13670
rect 29184 13456 29236 13462
rect 29184 13398 29236 13404
rect 29052 13268 29132 13274
rect 29000 13262 29132 13268
rect 29012 13246 29132 13262
rect 29012 12986 29040 13246
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 28908 12844 28960 12850
rect 28908 12786 28960 12792
rect 28397 12540 28705 12549
rect 28397 12538 28403 12540
rect 28459 12538 28483 12540
rect 28539 12538 28563 12540
rect 28619 12538 28643 12540
rect 28699 12538 28705 12540
rect 28459 12486 28461 12538
rect 28641 12486 28643 12538
rect 28397 12484 28403 12486
rect 28459 12484 28483 12486
rect 28539 12484 28563 12486
rect 28619 12484 28643 12486
rect 28699 12484 28705 12486
rect 28397 12475 28705 12484
rect 28092 12406 28304 12434
rect 28080 12096 28132 12102
rect 28080 12038 28132 12044
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 28092 11762 28120 12038
rect 28184 11898 28212 12038
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27988 11756 28040 11762
rect 27988 11698 28040 11704
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27356 10674 27384 11494
rect 27436 11280 27488 11286
rect 27436 11222 27488 11228
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27448 10062 27476 11222
rect 27540 11082 27568 11630
rect 27632 11218 27660 11698
rect 27804 11620 27856 11626
rect 27804 11562 27856 11568
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27632 11014 27660 11154
rect 27816 11150 27844 11562
rect 28276 11234 28304 12406
rect 28724 11620 28776 11626
rect 28724 11562 28776 11568
rect 28397 11452 28705 11461
rect 28397 11450 28403 11452
rect 28459 11450 28483 11452
rect 28539 11450 28563 11452
rect 28619 11450 28643 11452
rect 28699 11450 28705 11452
rect 28459 11398 28461 11450
rect 28641 11398 28643 11450
rect 28397 11396 28403 11398
rect 28459 11396 28483 11398
rect 28539 11396 28563 11398
rect 28619 11396 28643 11398
rect 28699 11396 28705 11398
rect 28397 11387 28705 11396
rect 28736 11268 28764 11562
rect 28184 11206 28304 11234
rect 28644 11240 28764 11268
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27816 11014 27844 11086
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27804 11008 27856 11014
rect 27804 10950 27856 10956
rect 27632 10554 27660 10950
rect 27632 10526 27752 10554
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27632 10266 27660 10406
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27724 10146 27752 10526
rect 27632 10118 27752 10146
rect 27816 10130 27844 10950
rect 28000 10810 28028 11086
rect 27988 10804 28040 10810
rect 27988 10746 28040 10752
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 27804 10124 27856 10130
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27632 9926 27660 10118
rect 27804 10066 27856 10072
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 26700 9648 26752 9654
rect 26700 9590 26752 9596
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26148 9104 26200 9110
rect 26148 9046 26200 9052
rect 26252 8974 26280 9318
rect 26620 9178 26648 9590
rect 27632 9586 27660 9862
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24320 7546 24348 8026
rect 24780 7886 24808 8230
rect 25240 7886 25268 8774
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25424 8090 25452 8434
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 26804 7886 26832 9318
rect 26974 9072 27030 9081
rect 26974 9007 27030 9016
rect 26988 8974 27016 9007
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 27632 8634 27660 9522
rect 27724 9042 27752 9998
rect 27816 9382 27844 10066
rect 27908 9722 27936 10610
rect 28000 10606 28028 10746
rect 27988 10600 28040 10606
rect 27988 10542 28040 10548
rect 27988 10192 28040 10198
rect 27988 10134 28040 10140
rect 28000 9926 28028 10134
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 28184 9586 28212 11206
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28276 10062 28304 11018
rect 28644 10606 28672 11240
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 28736 10674 28764 10950
rect 28816 10804 28868 10810
rect 28816 10746 28868 10752
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28632 10600 28684 10606
rect 28684 10548 28764 10554
rect 28632 10542 28764 10548
rect 28644 10526 28764 10542
rect 28397 10364 28705 10373
rect 28397 10362 28403 10364
rect 28459 10362 28483 10364
rect 28539 10362 28563 10364
rect 28619 10362 28643 10364
rect 28699 10362 28705 10364
rect 28459 10310 28461 10362
rect 28641 10310 28643 10362
rect 28397 10308 28403 10310
rect 28459 10308 28483 10310
rect 28539 10308 28563 10310
rect 28619 10308 28643 10310
rect 28699 10308 28705 10310
rect 28397 10299 28705 10308
rect 28736 10062 28764 10526
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27816 8974 27844 9318
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 27264 8090 27292 8434
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 27632 7886 27660 8570
rect 27816 8294 27844 8910
rect 27908 8838 27936 9318
rect 28397 9276 28705 9285
rect 28397 9274 28403 9276
rect 28459 9274 28483 9276
rect 28539 9274 28563 9276
rect 28619 9274 28643 9276
rect 28699 9274 28705 9276
rect 28459 9222 28461 9274
rect 28641 9222 28643 9274
rect 28397 9220 28403 9222
rect 28459 9220 28483 9222
rect 28539 9220 28563 9222
rect 28619 9220 28643 9222
rect 28699 9220 28705 9222
rect 28397 9211 28705 9220
rect 28172 9036 28224 9042
rect 28172 8978 28224 8984
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27816 7954 27844 8230
rect 28184 8090 28212 8978
rect 28736 8974 28764 9998
rect 28828 9586 28856 10746
rect 28920 10674 28948 12786
rect 29012 12782 29040 12922
rect 29196 12918 29224 13398
rect 29184 12912 29236 12918
rect 29184 12854 29236 12860
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 29000 12096 29052 12102
rect 29000 12038 29052 12044
rect 29012 11218 29040 12038
rect 29104 11626 29132 12174
rect 29276 12164 29328 12170
rect 29276 12106 29328 12112
rect 29092 11620 29144 11626
rect 29092 11562 29144 11568
rect 29000 11212 29052 11218
rect 29000 11154 29052 11160
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29196 10742 29224 11086
rect 29288 11082 29316 12106
rect 29380 11898 29408 13874
rect 29564 13530 29592 14894
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29656 13870 29684 14758
rect 29748 14278 29776 15098
rect 29828 14816 29880 14822
rect 29828 14758 29880 14764
rect 29840 14414 29868 14758
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29736 14272 29788 14278
rect 29736 14214 29788 14220
rect 29748 13938 29776 14214
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 29748 13410 29776 13874
rect 29460 13388 29512 13394
rect 29460 13330 29512 13336
rect 29656 13382 29776 13410
rect 29472 12306 29500 13330
rect 29656 13190 29684 13382
rect 29932 13326 29960 17478
rect 30024 17202 30052 17478
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 30300 17134 30328 17614
rect 30392 17270 30420 18022
rect 31116 17876 31168 17882
rect 31116 17818 31168 17824
rect 30380 17264 30432 17270
rect 30380 17206 30432 17212
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30472 16992 30524 16998
rect 30286 16960 30342 16969
rect 30342 16918 30420 16946
rect 30472 16934 30524 16940
rect 30286 16895 30342 16904
rect 30392 16182 30420 16918
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 30380 15632 30432 15638
rect 30208 15580 30380 15586
rect 30208 15574 30432 15580
rect 30208 15570 30420 15574
rect 30196 15564 30420 15570
rect 30248 15558 30420 15564
rect 30196 15506 30248 15512
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30024 15094 30052 15438
rect 30104 15428 30156 15434
rect 30104 15370 30156 15376
rect 30012 15088 30064 15094
rect 30012 15030 30064 15036
rect 30116 14346 30144 15370
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30104 14340 30156 14346
rect 30104 14282 30156 14288
rect 30392 13734 30420 15302
rect 30484 15026 30512 16934
rect 31128 16794 31156 17818
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 31036 15706 31064 16050
rect 31116 16040 31168 16046
rect 31116 15982 31168 15988
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 31128 15094 31156 15982
rect 31116 15088 31168 15094
rect 31116 15030 31168 15036
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 31128 14618 31156 15030
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 30472 14000 30524 14006
rect 30472 13942 30524 13948
rect 30380 13728 30432 13734
rect 30380 13670 30432 13676
rect 30012 13456 30064 13462
rect 30012 13398 30064 13404
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29656 12850 29684 13126
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 29840 12374 29868 12786
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29828 12368 29880 12374
rect 29828 12310 29880 12316
rect 29460 12300 29512 12306
rect 29460 12242 29512 12248
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29368 11892 29420 11898
rect 29368 11834 29420 11840
rect 29656 11762 29684 12174
rect 29736 12096 29788 12102
rect 29736 12038 29788 12044
rect 29748 11830 29776 12038
rect 29736 11824 29788 11830
rect 29736 11766 29788 11772
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29276 11076 29328 11082
rect 29276 11018 29328 11024
rect 29184 10736 29236 10742
rect 29184 10678 29236 10684
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 28816 9580 28868 9586
rect 28816 9522 28868 9528
rect 28920 8974 28948 10610
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 29012 9178 29040 10542
rect 29288 10538 29316 11018
rect 29276 10532 29328 10538
rect 29276 10474 29328 10480
rect 29656 10470 29684 11698
rect 29736 10668 29788 10674
rect 29840 10656 29868 12310
rect 29932 11694 29960 12582
rect 30024 12306 30052 13398
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30208 11898 30236 12174
rect 30196 11892 30248 11898
rect 30196 11834 30248 11840
rect 29920 11688 29972 11694
rect 29920 11630 29972 11636
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30208 11354 30236 11630
rect 30196 11348 30248 11354
rect 30196 11290 30248 11296
rect 30104 10736 30156 10742
rect 30104 10678 30156 10684
rect 29788 10628 29868 10656
rect 30012 10668 30064 10674
rect 29736 10610 29788 10616
rect 30012 10610 30064 10616
rect 29748 10470 29776 10610
rect 29644 10464 29696 10470
rect 29644 10406 29696 10412
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29472 9722 29500 10066
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29472 9586 29500 9658
rect 29460 9580 29512 9586
rect 29460 9522 29512 9528
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 29656 9042 29684 10406
rect 29748 9518 29776 10406
rect 30024 10130 30052 10610
rect 30012 10124 30064 10130
rect 30012 10066 30064 10072
rect 30116 10062 30144 10678
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30300 9586 30328 12718
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30392 11082 30420 12106
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30484 10554 30512 13942
rect 31404 13870 31432 14962
rect 31392 13864 31444 13870
rect 31392 13806 31444 13812
rect 30932 13524 30984 13530
rect 30932 13466 30984 13472
rect 30564 12844 30616 12850
rect 30564 12786 30616 12792
rect 30576 12442 30604 12786
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30760 11354 30788 12174
rect 30944 11354 30972 13466
rect 31024 11552 31076 11558
rect 31024 11494 31076 11500
rect 30748 11348 30800 11354
rect 30748 11290 30800 11296
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 30748 11076 30800 11082
rect 30748 11018 30800 11024
rect 30760 10674 30788 11018
rect 30748 10668 30800 10674
rect 30748 10610 30800 10616
rect 30564 10600 30616 10606
rect 30484 10548 30564 10554
rect 30484 10542 30616 10548
rect 30484 10526 30604 10542
rect 30484 9722 30512 10526
rect 30944 10130 30972 11290
rect 31036 11218 31064 11494
rect 31024 11212 31076 11218
rect 31024 11154 31076 11160
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 31036 10266 31064 10406
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 31128 10062 31156 10746
rect 31312 10674 31340 11086
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 30472 9716 30524 9722
rect 30472 9658 30524 9664
rect 30852 9654 30880 9930
rect 31128 9722 31156 9998
rect 31116 9716 31168 9722
rect 31116 9658 31168 9664
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 29736 9512 29788 9518
rect 29788 9460 29868 9466
rect 29736 9454 29868 9460
rect 29748 9438 29868 9454
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 29748 8974 29776 9318
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28908 8968 28960 8974
rect 28908 8910 28960 8916
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29840 8634 29868 9438
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 30300 8566 30328 9522
rect 31496 9382 31524 19450
rect 31588 18766 31616 19654
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31680 18358 31708 20198
rect 31668 18352 31720 18358
rect 31668 18294 31720 18300
rect 31576 18080 31628 18086
rect 31576 18022 31628 18028
rect 31588 17610 31616 18022
rect 31758 17912 31814 17921
rect 31758 17847 31814 17856
rect 31576 17604 31628 17610
rect 31576 17546 31628 17552
rect 31668 16448 31720 16454
rect 31668 16390 31720 16396
rect 31680 15366 31708 16390
rect 31668 15360 31720 15366
rect 31668 15302 31720 15308
rect 31772 14074 31800 17847
rect 31864 17678 31892 21406
rect 32318 20700 32626 20709
rect 32318 20698 32324 20700
rect 32380 20698 32404 20700
rect 32460 20698 32484 20700
rect 32540 20698 32564 20700
rect 32620 20698 32626 20700
rect 32380 20646 32382 20698
rect 32562 20646 32564 20698
rect 32318 20644 32324 20646
rect 32380 20644 32404 20646
rect 32460 20644 32484 20646
rect 32540 20644 32564 20646
rect 32620 20644 32626 20646
rect 32318 20635 32626 20644
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31852 17672 31904 17678
rect 31852 17614 31904 17620
rect 31852 17536 31904 17542
rect 31852 17478 31904 17484
rect 31864 16590 31892 17478
rect 31852 16584 31904 16590
rect 31852 16526 31904 16532
rect 31956 16250 31984 19790
rect 32318 19612 32626 19621
rect 32318 19610 32324 19612
rect 32380 19610 32404 19612
rect 32460 19610 32484 19612
rect 32540 19610 32564 19612
rect 32620 19610 32626 19612
rect 32380 19558 32382 19610
rect 32562 19558 32564 19610
rect 32318 19556 32324 19558
rect 32380 19556 32404 19558
rect 32460 19556 32484 19558
rect 32540 19556 32564 19558
rect 32620 19556 32626 19558
rect 32318 19547 32626 19556
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 31944 16244 31996 16250
rect 31944 16186 31996 16192
rect 31760 14068 31812 14074
rect 31760 14010 31812 14016
rect 32048 12918 32076 18566
rect 32318 18524 32626 18533
rect 32318 18522 32324 18524
rect 32380 18522 32404 18524
rect 32460 18522 32484 18524
rect 32540 18522 32564 18524
rect 32620 18522 32626 18524
rect 32380 18470 32382 18522
rect 32562 18470 32564 18522
rect 32318 18468 32324 18470
rect 32380 18468 32404 18470
rect 32460 18468 32484 18470
rect 32540 18468 32564 18470
rect 32620 18468 32626 18470
rect 32318 18459 32626 18468
rect 32318 17436 32626 17445
rect 32318 17434 32324 17436
rect 32380 17434 32404 17436
rect 32460 17434 32484 17436
rect 32540 17434 32564 17436
rect 32620 17434 32626 17436
rect 32380 17382 32382 17434
rect 32562 17382 32564 17434
rect 32318 17380 32324 17382
rect 32380 17380 32404 17382
rect 32460 17380 32484 17382
rect 32540 17380 32564 17382
rect 32620 17380 32626 17382
rect 32318 17371 32626 17380
rect 32318 16348 32626 16357
rect 32318 16346 32324 16348
rect 32380 16346 32404 16348
rect 32460 16346 32484 16348
rect 32540 16346 32564 16348
rect 32620 16346 32626 16348
rect 32380 16294 32382 16346
rect 32562 16294 32564 16346
rect 32318 16292 32324 16294
rect 32380 16292 32404 16294
rect 32460 16292 32484 16294
rect 32540 16292 32564 16294
rect 32620 16292 32626 16294
rect 32318 16283 32626 16292
rect 32318 15260 32626 15269
rect 32318 15258 32324 15260
rect 32380 15258 32404 15260
rect 32460 15258 32484 15260
rect 32540 15258 32564 15260
rect 32620 15258 32626 15260
rect 32380 15206 32382 15258
rect 32562 15206 32564 15258
rect 32318 15204 32324 15206
rect 32380 15204 32404 15206
rect 32460 15204 32484 15206
rect 32540 15204 32564 15206
rect 32620 15204 32626 15206
rect 32318 15195 32626 15204
rect 32318 14172 32626 14181
rect 32318 14170 32324 14172
rect 32380 14170 32404 14172
rect 32460 14170 32484 14172
rect 32540 14170 32564 14172
rect 32620 14170 32626 14172
rect 32380 14118 32382 14170
rect 32562 14118 32564 14170
rect 32318 14116 32324 14118
rect 32380 14116 32404 14118
rect 32460 14116 32484 14118
rect 32540 14116 32564 14118
rect 32620 14116 32626 14118
rect 32318 14107 32626 14116
rect 32318 13084 32626 13093
rect 32318 13082 32324 13084
rect 32380 13082 32404 13084
rect 32460 13082 32484 13084
rect 32540 13082 32564 13084
rect 32620 13082 32626 13084
rect 32380 13030 32382 13082
rect 32562 13030 32564 13082
rect 32318 13028 32324 13030
rect 32380 13028 32404 13030
rect 32460 13028 32484 13030
rect 32540 13028 32564 13030
rect 32620 13028 32626 13030
rect 32318 13019 32626 13028
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 32318 11996 32626 12005
rect 32318 11994 32324 11996
rect 32380 11994 32404 11996
rect 32460 11994 32484 11996
rect 32540 11994 32564 11996
rect 32620 11994 32626 11996
rect 32380 11942 32382 11994
rect 32562 11942 32564 11994
rect 32318 11940 32324 11942
rect 32380 11940 32404 11942
rect 32460 11940 32484 11942
rect 32540 11940 32564 11942
rect 32620 11940 32626 11942
rect 32318 11931 32626 11940
rect 31944 11280 31996 11286
rect 31944 11222 31996 11228
rect 31760 10668 31812 10674
rect 31760 10610 31812 10616
rect 31772 10266 31800 10610
rect 31760 10260 31812 10266
rect 31760 10202 31812 10208
rect 31956 10062 31984 11222
rect 32318 10908 32626 10917
rect 32318 10906 32324 10908
rect 32380 10906 32404 10908
rect 32460 10906 32484 10908
rect 32540 10906 32564 10908
rect 32620 10906 32626 10908
rect 32380 10854 32382 10906
rect 32562 10854 32564 10906
rect 32318 10852 32324 10854
rect 32380 10852 32404 10854
rect 32460 10852 32484 10854
rect 32540 10852 32564 10854
rect 32620 10852 32626 10854
rect 32318 10843 32626 10852
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 32318 9820 32626 9829
rect 32318 9818 32324 9820
rect 32380 9818 32404 9820
rect 32460 9818 32484 9820
rect 32540 9818 32564 9820
rect 32620 9818 32626 9820
rect 32380 9766 32382 9818
rect 32562 9766 32564 9818
rect 32318 9764 32324 9766
rect 32380 9764 32404 9766
rect 32460 9764 32484 9766
rect 32540 9764 32564 9766
rect 32620 9764 32626 9766
rect 32318 9755 32626 9764
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30288 8560 30340 8566
rect 30288 8502 30340 8508
rect 30392 8498 30420 8774
rect 32318 8732 32626 8741
rect 32318 8730 32324 8732
rect 32380 8730 32404 8732
rect 32460 8730 32484 8732
rect 32540 8730 32564 8732
rect 32620 8730 32626 8732
rect 32380 8678 32382 8730
rect 32562 8678 32564 8730
rect 32318 8676 32324 8678
rect 32380 8676 32404 8678
rect 32460 8676 32484 8678
rect 32540 8676 32564 8678
rect 32620 8676 32626 8678
rect 32318 8667 32626 8676
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 28397 8188 28705 8197
rect 28397 8186 28403 8188
rect 28459 8186 28483 8188
rect 28539 8186 28563 8188
rect 28619 8186 28643 8188
rect 28699 8186 28705 8188
rect 28459 8134 28461 8186
rect 28641 8134 28643 8186
rect 28397 8132 28403 8134
rect 28459 8132 28483 8134
rect 28539 8132 28563 8134
rect 28619 8132 28643 8134
rect 28699 8132 28705 8134
rect 28397 8123 28705 8132
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24412 7546 24440 7686
rect 24476 7644 24784 7653
rect 24476 7642 24482 7644
rect 24538 7642 24562 7644
rect 24618 7642 24642 7644
rect 24698 7642 24722 7644
rect 24778 7642 24784 7644
rect 24538 7590 24540 7642
rect 24720 7590 24722 7642
rect 24476 7588 24482 7590
rect 24538 7588 24562 7590
rect 24618 7588 24642 7590
rect 24698 7588 24722 7590
rect 24778 7588 24784 7590
rect 24476 7579 24784 7588
rect 32318 7644 32626 7653
rect 32318 7642 32324 7644
rect 32380 7642 32404 7644
rect 32460 7642 32484 7644
rect 32540 7642 32564 7644
rect 32620 7642 32626 7644
rect 32380 7590 32382 7642
rect 32562 7590 32564 7642
rect 32318 7588 32324 7590
rect 32380 7588 32404 7590
rect 32460 7588 32484 7590
rect 32540 7588 32564 7590
rect 32620 7588 32626 7590
rect 32318 7579 32626 7588
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24596 7410 24900 7426
rect 24584 7404 24912 7410
rect 24636 7398 24860 7404
rect 24584 7346 24636 7352
rect 24860 7346 24912 7352
rect 24596 7274 24624 7346
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 24584 7268 24636 7274
rect 24584 7210 24636 7216
rect 24676 7268 24728 7274
rect 24676 7210 24728 7216
rect 24688 7002 24716 7210
rect 28397 7100 28705 7109
rect 28397 7098 28403 7100
rect 28459 7098 28483 7100
rect 28539 7098 28563 7100
rect 28619 7098 28643 7100
rect 28699 7098 28705 7100
rect 28459 7046 28461 7098
rect 28641 7046 28643 7098
rect 28397 7044 28403 7046
rect 28459 7044 28483 7046
rect 28539 7044 28563 7046
rect 28619 7044 28643 7046
rect 28699 7044 28705 7046
rect 28397 7035 28705 7044
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 24476 6556 24784 6565
rect 24476 6554 24482 6556
rect 24538 6554 24562 6556
rect 24618 6554 24642 6556
rect 24698 6554 24722 6556
rect 24778 6554 24784 6556
rect 24538 6502 24540 6554
rect 24720 6502 24722 6554
rect 24476 6500 24482 6502
rect 24538 6500 24562 6502
rect 24618 6500 24642 6502
rect 24698 6500 24722 6502
rect 24778 6500 24784 6502
rect 24476 6491 24784 6500
rect 32318 6556 32626 6565
rect 32318 6554 32324 6556
rect 32380 6554 32404 6556
rect 32460 6554 32484 6556
rect 32540 6554 32564 6556
rect 32620 6554 32626 6556
rect 32380 6502 32382 6554
rect 32562 6502 32564 6554
rect 32318 6500 32324 6502
rect 32380 6500 32404 6502
rect 32460 6500 32484 6502
rect 32540 6500 32564 6502
rect 32620 6500 32626 6502
rect 32318 6491 32626 6500
rect 28397 6012 28705 6021
rect 28397 6010 28403 6012
rect 28459 6010 28483 6012
rect 28539 6010 28563 6012
rect 28619 6010 28643 6012
rect 28699 6010 28705 6012
rect 28459 5958 28461 6010
rect 28641 5958 28643 6010
rect 28397 5956 28403 5958
rect 28459 5956 28483 5958
rect 28539 5956 28563 5958
rect 28619 5956 28643 5958
rect 28699 5956 28705 5958
rect 28397 5947 28705 5956
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21744 5302 21772 5510
rect 21836 5370 21864 5646
rect 24476 5468 24784 5477
rect 24476 5466 24482 5468
rect 24538 5466 24562 5468
rect 24618 5466 24642 5468
rect 24698 5466 24722 5468
rect 24778 5466 24784 5468
rect 24538 5414 24540 5466
rect 24720 5414 24722 5466
rect 24476 5412 24482 5414
rect 24538 5412 24562 5414
rect 24618 5412 24642 5414
rect 24698 5412 24722 5414
rect 24778 5412 24784 5414
rect 24476 5403 24784 5412
rect 32318 5468 32626 5477
rect 32318 5466 32324 5468
rect 32380 5466 32404 5468
rect 32460 5466 32484 5468
rect 32540 5466 32564 5468
rect 32620 5466 32626 5468
rect 32380 5414 32382 5466
rect 32562 5414 32564 5466
rect 32318 5412 32324 5414
rect 32380 5412 32404 5414
rect 32460 5412 32484 5414
rect 32540 5412 32564 5414
rect 32620 5412 32626 5414
rect 32318 5403 32626 5412
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 4871 4924 5179 4933
rect 4871 4922 4877 4924
rect 4933 4922 4957 4924
rect 5013 4922 5037 4924
rect 5093 4922 5117 4924
rect 5173 4922 5179 4924
rect 4933 4870 4935 4922
rect 5115 4870 5117 4922
rect 4871 4868 4877 4870
rect 4933 4868 4957 4870
rect 5013 4868 5037 4870
rect 5093 4868 5117 4870
rect 5173 4868 5179 4870
rect 4871 4859 5179 4868
rect 12713 4924 13021 4933
rect 12713 4922 12719 4924
rect 12775 4922 12799 4924
rect 12855 4922 12879 4924
rect 12935 4922 12959 4924
rect 13015 4922 13021 4924
rect 12775 4870 12777 4922
rect 12957 4870 12959 4922
rect 12713 4868 12719 4870
rect 12775 4868 12799 4870
rect 12855 4868 12879 4870
rect 12935 4868 12959 4870
rect 13015 4868 13021 4870
rect 12713 4859 13021 4868
rect 20555 4924 20863 4933
rect 20555 4922 20561 4924
rect 20617 4922 20641 4924
rect 20697 4922 20721 4924
rect 20777 4922 20801 4924
rect 20857 4922 20863 4924
rect 20617 4870 20619 4922
rect 20799 4870 20801 4922
rect 20555 4868 20561 4870
rect 20617 4868 20641 4870
rect 20697 4868 20721 4870
rect 20777 4868 20801 4870
rect 20857 4868 20863 4870
rect 20555 4859 20863 4868
rect 28397 4924 28705 4933
rect 28397 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28643 4924
rect 28699 4922 28705 4924
rect 28459 4870 28461 4922
rect 28641 4870 28643 4922
rect 28397 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28643 4870
rect 28699 4868 28705 4870
rect 28397 4859 28705 4868
rect 8792 4380 9100 4389
rect 8792 4378 8798 4380
rect 8854 4378 8878 4380
rect 8934 4378 8958 4380
rect 9014 4378 9038 4380
rect 9094 4378 9100 4380
rect 8854 4326 8856 4378
rect 9036 4326 9038 4378
rect 8792 4324 8798 4326
rect 8854 4324 8878 4326
rect 8934 4324 8958 4326
rect 9014 4324 9038 4326
rect 9094 4324 9100 4326
rect 8792 4315 9100 4324
rect 16634 4380 16942 4389
rect 16634 4378 16640 4380
rect 16696 4378 16720 4380
rect 16776 4378 16800 4380
rect 16856 4378 16880 4380
rect 16936 4378 16942 4380
rect 16696 4326 16698 4378
rect 16878 4326 16880 4378
rect 16634 4324 16640 4326
rect 16696 4324 16720 4326
rect 16776 4324 16800 4326
rect 16856 4324 16880 4326
rect 16936 4324 16942 4326
rect 16634 4315 16942 4324
rect 24476 4380 24784 4389
rect 24476 4378 24482 4380
rect 24538 4378 24562 4380
rect 24618 4378 24642 4380
rect 24698 4378 24722 4380
rect 24778 4378 24784 4380
rect 24538 4326 24540 4378
rect 24720 4326 24722 4378
rect 24476 4324 24482 4326
rect 24538 4324 24562 4326
rect 24618 4324 24642 4326
rect 24698 4324 24722 4326
rect 24778 4324 24784 4326
rect 24476 4315 24784 4324
rect 32318 4380 32626 4389
rect 32318 4378 32324 4380
rect 32380 4378 32404 4380
rect 32460 4378 32484 4380
rect 32540 4378 32564 4380
rect 32620 4378 32626 4380
rect 32380 4326 32382 4378
rect 32562 4326 32564 4378
rect 32318 4324 32324 4326
rect 32380 4324 32404 4326
rect 32460 4324 32484 4326
rect 32540 4324 32564 4326
rect 32620 4324 32626 4326
rect 32318 4315 32626 4324
rect 4871 3836 5179 3845
rect 4871 3834 4877 3836
rect 4933 3834 4957 3836
rect 5013 3834 5037 3836
rect 5093 3834 5117 3836
rect 5173 3834 5179 3836
rect 4933 3782 4935 3834
rect 5115 3782 5117 3834
rect 4871 3780 4877 3782
rect 4933 3780 4957 3782
rect 5013 3780 5037 3782
rect 5093 3780 5117 3782
rect 5173 3780 5179 3782
rect 4871 3771 5179 3780
rect 12713 3836 13021 3845
rect 12713 3834 12719 3836
rect 12775 3834 12799 3836
rect 12855 3834 12879 3836
rect 12935 3834 12959 3836
rect 13015 3834 13021 3836
rect 12775 3782 12777 3834
rect 12957 3782 12959 3834
rect 12713 3780 12719 3782
rect 12775 3780 12799 3782
rect 12855 3780 12879 3782
rect 12935 3780 12959 3782
rect 13015 3780 13021 3782
rect 12713 3771 13021 3780
rect 20555 3836 20863 3845
rect 20555 3834 20561 3836
rect 20617 3834 20641 3836
rect 20697 3834 20721 3836
rect 20777 3834 20801 3836
rect 20857 3834 20863 3836
rect 20617 3782 20619 3834
rect 20799 3782 20801 3834
rect 20555 3780 20561 3782
rect 20617 3780 20641 3782
rect 20697 3780 20721 3782
rect 20777 3780 20801 3782
rect 20857 3780 20863 3782
rect 20555 3771 20863 3780
rect 28397 3836 28705 3845
rect 28397 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28643 3836
rect 28699 3834 28705 3836
rect 28459 3782 28461 3834
rect 28641 3782 28643 3834
rect 28397 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28643 3782
rect 28699 3780 28705 3782
rect 28397 3771 28705 3780
rect 8792 3292 9100 3301
rect 8792 3290 8798 3292
rect 8854 3290 8878 3292
rect 8934 3290 8958 3292
rect 9014 3290 9038 3292
rect 9094 3290 9100 3292
rect 8854 3238 8856 3290
rect 9036 3238 9038 3290
rect 8792 3236 8798 3238
rect 8854 3236 8878 3238
rect 8934 3236 8958 3238
rect 9014 3236 9038 3238
rect 9094 3236 9100 3238
rect 8792 3227 9100 3236
rect 16634 3292 16942 3301
rect 16634 3290 16640 3292
rect 16696 3290 16720 3292
rect 16776 3290 16800 3292
rect 16856 3290 16880 3292
rect 16936 3290 16942 3292
rect 16696 3238 16698 3290
rect 16878 3238 16880 3290
rect 16634 3236 16640 3238
rect 16696 3236 16720 3238
rect 16776 3236 16800 3238
rect 16856 3236 16880 3238
rect 16936 3236 16942 3238
rect 16634 3227 16942 3236
rect 24476 3292 24784 3301
rect 24476 3290 24482 3292
rect 24538 3290 24562 3292
rect 24618 3290 24642 3292
rect 24698 3290 24722 3292
rect 24778 3290 24784 3292
rect 24538 3238 24540 3290
rect 24720 3238 24722 3290
rect 24476 3236 24482 3238
rect 24538 3236 24562 3238
rect 24618 3236 24642 3238
rect 24698 3236 24722 3238
rect 24778 3236 24784 3238
rect 24476 3227 24784 3236
rect 32318 3292 32626 3301
rect 32318 3290 32324 3292
rect 32380 3290 32404 3292
rect 32460 3290 32484 3292
rect 32540 3290 32564 3292
rect 32620 3290 32626 3292
rect 32380 3238 32382 3290
rect 32562 3238 32564 3290
rect 32318 3236 32324 3238
rect 32380 3236 32404 3238
rect 32460 3236 32484 3238
rect 32540 3236 32564 3238
rect 32620 3236 32626 3238
rect 32318 3227 32626 3236
rect 4871 2748 5179 2757
rect 4871 2746 4877 2748
rect 4933 2746 4957 2748
rect 5013 2746 5037 2748
rect 5093 2746 5117 2748
rect 5173 2746 5179 2748
rect 4933 2694 4935 2746
rect 5115 2694 5117 2746
rect 4871 2692 4877 2694
rect 4933 2692 4957 2694
rect 5013 2692 5037 2694
rect 5093 2692 5117 2694
rect 5173 2692 5179 2694
rect 4871 2683 5179 2692
rect 12713 2748 13021 2757
rect 12713 2746 12719 2748
rect 12775 2746 12799 2748
rect 12855 2746 12879 2748
rect 12935 2746 12959 2748
rect 13015 2746 13021 2748
rect 12775 2694 12777 2746
rect 12957 2694 12959 2746
rect 12713 2692 12719 2694
rect 12775 2692 12799 2694
rect 12855 2692 12879 2694
rect 12935 2692 12959 2694
rect 13015 2692 13021 2694
rect 12713 2683 13021 2692
rect 20555 2748 20863 2757
rect 20555 2746 20561 2748
rect 20617 2746 20641 2748
rect 20697 2746 20721 2748
rect 20777 2746 20801 2748
rect 20857 2746 20863 2748
rect 20617 2694 20619 2746
rect 20799 2694 20801 2746
rect 20555 2692 20561 2694
rect 20617 2692 20641 2694
rect 20697 2692 20721 2694
rect 20777 2692 20801 2694
rect 20857 2692 20863 2694
rect 20555 2683 20863 2692
rect 28397 2748 28705 2757
rect 28397 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28643 2748
rect 28699 2746 28705 2748
rect 28459 2694 28461 2746
rect 28641 2694 28643 2746
rect 28397 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28643 2694
rect 28699 2692 28705 2694
rect 28397 2683 28705 2692
rect 8792 2204 9100 2213
rect 8792 2202 8798 2204
rect 8854 2202 8878 2204
rect 8934 2202 8958 2204
rect 9014 2202 9038 2204
rect 9094 2202 9100 2204
rect 8854 2150 8856 2202
rect 9036 2150 9038 2202
rect 8792 2148 8798 2150
rect 8854 2148 8878 2150
rect 8934 2148 8958 2150
rect 9014 2148 9038 2150
rect 9094 2148 9100 2150
rect 8792 2139 9100 2148
rect 16634 2204 16942 2213
rect 16634 2202 16640 2204
rect 16696 2202 16720 2204
rect 16776 2202 16800 2204
rect 16856 2202 16880 2204
rect 16936 2202 16942 2204
rect 16696 2150 16698 2202
rect 16878 2150 16880 2202
rect 16634 2148 16640 2150
rect 16696 2148 16720 2150
rect 16776 2148 16800 2150
rect 16856 2148 16880 2150
rect 16936 2148 16942 2150
rect 16634 2139 16942 2148
rect 24476 2204 24784 2213
rect 24476 2202 24482 2204
rect 24538 2202 24562 2204
rect 24618 2202 24642 2204
rect 24698 2202 24722 2204
rect 24778 2202 24784 2204
rect 24538 2150 24540 2202
rect 24720 2150 24722 2202
rect 24476 2148 24482 2150
rect 24538 2148 24562 2150
rect 24618 2148 24642 2150
rect 24698 2148 24722 2150
rect 24778 2148 24784 2150
rect 24476 2139 24784 2148
rect 32318 2204 32626 2213
rect 32318 2202 32324 2204
rect 32380 2202 32404 2204
rect 32460 2202 32484 2204
rect 32540 2202 32564 2204
rect 32620 2202 32626 2204
rect 32380 2150 32382 2202
rect 32562 2150 32564 2202
rect 32318 2148 32324 2150
rect 32380 2148 32404 2150
rect 32460 2148 32484 2150
rect 32540 2148 32564 2150
rect 32620 2148 32626 2150
rect 32318 2139 32626 2148
rect 4871 1660 5179 1669
rect 4871 1658 4877 1660
rect 4933 1658 4957 1660
rect 5013 1658 5037 1660
rect 5093 1658 5117 1660
rect 5173 1658 5179 1660
rect 4933 1606 4935 1658
rect 5115 1606 5117 1658
rect 4871 1604 4877 1606
rect 4933 1604 4957 1606
rect 5013 1604 5037 1606
rect 5093 1604 5117 1606
rect 5173 1604 5179 1606
rect 4871 1595 5179 1604
rect 12713 1660 13021 1669
rect 12713 1658 12719 1660
rect 12775 1658 12799 1660
rect 12855 1658 12879 1660
rect 12935 1658 12959 1660
rect 13015 1658 13021 1660
rect 12775 1606 12777 1658
rect 12957 1606 12959 1658
rect 12713 1604 12719 1606
rect 12775 1604 12799 1606
rect 12855 1604 12879 1606
rect 12935 1604 12959 1606
rect 13015 1604 13021 1606
rect 12713 1595 13021 1604
rect 20555 1660 20863 1669
rect 20555 1658 20561 1660
rect 20617 1658 20641 1660
rect 20697 1658 20721 1660
rect 20777 1658 20801 1660
rect 20857 1658 20863 1660
rect 20617 1606 20619 1658
rect 20799 1606 20801 1658
rect 20555 1604 20561 1606
rect 20617 1604 20641 1606
rect 20697 1604 20721 1606
rect 20777 1604 20801 1606
rect 20857 1604 20863 1606
rect 20555 1595 20863 1604
rect 28397 1660 28705 1669
rect 28397 1658 28403 1660
rect 28459 1658 28483 1660
rect 28539 1658 28563 1660
rect 28619 1658 28643 1660
rect 28699 1658 28705 1660
rect 28459 1606 28461 1658
rect 28641 1606 28643 1658
rect 28397 1604 28403 1606
rect 28459 1604 28483 1606
rect 28539 1604 28563 1606
rect 28619 1604 28643 1606
rect 28699 1604 28705 1606
rect 28397 1595 28705 1604
rect 8792 1116 9100 1125
rect 8792 1114 8798 1116
rect 8854 1114 8878 1116
rect 8934 1114 8958 1116
rect 9014 1114 9038 1116
rect 9094 1114 9100 1116
rect 8854 1062 8856 1114
rect 9036 1062 9038 1114
rect 8792 1060 8798 1062
rect 8854 1060 8878 1062
rect 8934 1060 8958 1062
rect 9014 1060 9038 1062
rect 9094 1060 9100 1062
rect 8792 1051 9100 1060
rect 16634 1116 16942 1125
rect 16634 1114 16640 1116
rect 16696 1114 16720 1116
rect 16776 1114 16800 1116
rect 16856 1114 16880 1116
rect 16936 1114 16942 1116
rect 16696 1062 16698 1114
rect 16878 1062 16880 1114
rect 16634 1060 16640 1062
rect 16696 1060 16720 1062
rect 16776 1060 16800 1062
rect 16856 1060 16880 1062
rect 16936 1060 16942 1062
rect 16634 1051 16942 1060
rect 24476 1116 24784 1125
rect 24476 1114 24482 1116
rect 24538 1114 24562 1116
rect 24618 1114 24642 1116
rect 24698 1114 24722 1116
rect 24778 1114 24784 1116
rect 24538 1062 24540 1114
rect 24720 1062 24722 1114
rect 24476 1060 24482 1062
rect 24538 1060 24562 1062
rect 24618 1060 24642 1062
rect 24698 1060 24722 1062
rect 24778 1060 24784 1062
rect 24476 1051 24784 1060
rect 32318 1116 32626 1125
rect 32318 1114 32324 1116
rect 32380 1114 32404 1116
rect 32460 1114 32484 1116
rect 32540 1114 32564 1116
rect 32620 1114 32626 1116
rect 32380 1062 32382 1114
rect 32562 1062 32564 1114
rect 32318 1060 32324 1062
rect 32380 1060 32404 1062
rect 32460 1060 32484 1062
rect 32540 1060 32564 1062
rect 32620 1060 32626 1062
rect 32318 1051 32626 1060
<< via2 >>
rect 2962 21392 3018 21448
rect 4434 21392 4490 21448
rect 4802 21392 4858 21448
rect 5538 21392 5594 21448
rect 6090 21392 6146 21448
rect 8206 21392 8262 21448
rect 9678 21392 9734 21448
rect 11794 21392 11850 21448
rect 13818 21392 13874 21448
rect 14186 21392 14242 21448
rect 15842 21392 15898 21448
rect 28262 21392 28318 21448
rect 28722 21392 28778 21448
rect 29458 21392 29514 21448
rect 31666 21392 31722 21448
rect 4877 20154 4933 20156
rect 4957 20154 5013 20156
rect 5037 20154 5093 20156
rect 5117 20154 5173 20156
rect 4877 20102 4923 20154
rect 4923 20102 4933 20154
rect 4957 20102 4987 20154
rect 4987 20102 4999 20154
rect 4999 20102 5013 20154
rect 5037 20102 5051 20154
rect 5051 20102 5063 20154
rect 5063 20102 5093 20154
rect 5117 20102 5127 20154
rect 5127 20102 5173 20154
rect 4877 20100 4933 20102
rect 4957 20100 5013 20102
rect 5037 20100 5093 20102
rect 5117 20100 5173 20102
rect 1766 19508 1822 19544
rect 1766 19488 1768 19508
rect 1768 19488 1820 19508
rect 1820 19488 1822 19508
rect 1582 17856 1638 17912
rect 3514 17856 3570 17912
rect 4877 19066 4933 19068
rect 4957 19066 5013 19068
rect 5037 19066 5093 19068
rect 5117 19066 5173 19068
rect 4877 19014 4923 19066
rect 4923 19014 4933 19066
rect 4957 19014 4987 19066
rect 4987 19014 4999 19066
rect 4999 19014 5013 19066
rect 5037 19014 5051 19066
rect 5051 19014 5063 19066
rect 5063 19014 5093 19066
rect 5117 19014 5127 19066
rect 5127 19014 5173 19066
rect 4877 19012 4933 19014
rect 4957 19012 5013 19014
rect 5037 19012 5093 19014
rect 5117 19012 5173 19014
rect 8114 20596 8170 20632
rect 8114 20576 8116 20596
rect 8116 20576 8168 20596
rect 8168 20576 8170 20596
rect 9494 20848 9550 20904
rect 8798 20698 8854 20700
rect 8878 20698 8934 20700
rect 8958 20698 9014 20700
rect 9038 20698 9094 20700
rect 8798 20646 8844 20698
rect 8844 20646 8854 20698
rect 8878 20646 8908 20698
rect 8908 20646 8920 20698
rect 8920 20646 8934 20698
rect 8958 20646 8972 20698
rect 8972 20646 8984 20698
rect 8984 20646 9014 20698
rect 9038 20646 9048 20698
rect 9048 20646 9094 20698
rect 8798 20644 8854 20646
rect 8878 20644 8934 20646
rect 8958 20644 9014 20646
rect 9038 20644 9094 20646
rect 11058 21256 11114 21312
rect 11702 21256 11758 21312
rect 4877 17978 4933 17980
rect 4957 17978 5013 17980
rect 5037 17978 5093 17980
rect 5117 17978 5173 17980
rect 4877 17926 4923 17978
rect 4923 17926 4933 17978
rect 4957 17926 4987 17978
rect 4987 17926 4999 17978
rect 4999 17926 5013 17978
rect 5037 17926 5051 17978
rect 5051 17926 5063 17978
rect 5063 17926 5093 17978
rect 5117 17926 5127 17978
rect 5127 17926 5173 17978
rect 4877 17924 4933 17926
rect 4957 17924 5013 17926
rect 5037 17924 5093 17926
rect 5117 17924 5173 17926
rect 4877 16890 4933 16892
rect 4957 16890 5013 16892
rect 5037 16890 5093 16892
rect 5117 16890 5173 16892
rect 4877 16838 4923 16890
rect 4923 16838 4933 16890
rect 4957 16838 4987 16890
rect 4987 16838 4999 16890
rect 4999 16838 5013 16890
rect 5037 16838 5051 16890
rect 5051 16838 5063 16890
rect 5063 16838 5093 16890
rect 5117 16838 5127 16890
rect 5127 16838 5173 16890
rect 4877 16836 4933 16838
rect 4957 16836 5013 16838
rect 5037 16836 5093 16838
rect 5117 16836 5173 16838
rect 7102 17076 7104 17096
rect 7104 17076 7156 17096
rect 7156 17076 7158 17096
rect 7102 17040 7158 17076
rect 8798 19610 8854 19612
rect 8878 19610 8934 19612
rect 8958 19610 9014 19612
rect 9038 19610 9094 19612
rect 8798 19558 8844 19610
rect 8844 19558 8854 19610
rect 8878 19558 8908 19610
rect 8908 19558 8920 19610
rect 8920 19558 8934 19610
rect 8958 19558 8972 19610
rect 8972 19558 8984 19610
rect 8984 19558 9014 19610
rect 9038 19558 9048 19610
rect 9048 19558 9094 19610
rect 8798 19556 8854 19558
rect 8878 19556 8934 19558
rect 8958 19556 9014 19558
rect 9038 19556 9094 19558
rect 4877 15802 4933 15804
rect 4957 15802 5013 15804
rect 5037 15802 5093 15804
rect 5117 15802 5173 15804
rect 4877 15750 4923 15802
rect 4923 15750 4933 15802
rect 4957 15750 4987 15802
rect 4987 15750 4999 15802
rect 4999 15750 5013 15802
rect 5037 15750 5051 15802
rect 5051 15750 5063 15802
rect 5063 15750 5093 15802
rect 5117 15750 5127 15802
rect 5127 15750 5173 15802
rect 4877 15748 4933 15750
rect 4957 15748 5013 15750
rect 5037 15748 5093 15750
rect 5117 15748 5173 15750
rect 4877 14714 4933 14716
rect 4957 14714 5013 14716
rect 5037 14714 5093 14716
rect 5117 14714 5173 14716
rect 4877 14662 4923 14714
rect 4923 14662 4933 14714
rect 4957 14662 4987 14714
rect 4987 14662 4999 14714
rect 4999 14662 5013 14714
rect 5037 14662 5051 14714
rect 5051 14662 5063 14714
rect 5063 14662 5093 14714
rect 5117 14662 5127 14714
rect 5127 14662 5173 14714
rect 4877 14660 4933 14662
rect 4957 14660 5013 14662
rect 5037 14660 5093 14662
rect 5117 14660 5173 14662
rect 4877 13626 4933 13628
rect 4957 13626 5013 13628
rect 5037 13626 5093 13628
rect 5117 13626 5173 13628
rect 4877 13574 4923 13626
rect 4923 13574 4933 13626
rect 4957 13574 4987 13626
rect 4987 13574 4999 13626
rect 4999 13574 5013 13626
rect 5037 13574 5051 13626
rect 5051 13574 5063 13626
rect 5063 13574 5093 13626
rect 5117 13574 5127 13626
rect 5127 13574 5173 13626
rect 4877 13572 4933 13574
rect 4957 13572 5013 13574
rect 5037 13572 5093 13574
rect 5117 13572 5173 13574
rect 4877 12538 4933 12540
rect 4957 12538 5013 12540
rect 5037 12538 5093 12540
rect 5117 12538 5173 12540
rect 4877 12486 4923 12538
rect 4923 12486 4933 12538
rect 4957 12486 4987 12538
rect 4987 12486 4999 12538
rect 4999 12486 5013 12538
rect 5037 12486 5051 12538
rect 5051 12486 5063 12538
rect 5063 12486 5093 12538
rect 5117 12486 5127 12538
rect 5127 12486 5173 12538
rect 4877 12484 4933 12486
rect 4957 12484 5013 12486
rect 5037 12484 5093 12486
rect 5117 12484 5173 12486
rect 4877 11450 4933 11452
rect 4957 11450 5013 11452
rect 5037 11450 5093 11452
rect 5117 11450 5173 11452
rect 4877 11398 4923 11450
rect 4923 11398 4933 11450
rect 4957 11398 4987 11450
rect 4987 11398 4999 11450
rect 4999 11398 5013 11450
rect 5037 11398 5051 11450
rect 5051 11398 5063 11450
rect 5063 11398 5093 11450
rect 5117 11398 5127 11450
rect 5127 11398 5173 11450
rect 4877 11396 4933 11398
rect 4957 11396 5013 11398
rect 5037 11396 5093 11398
rect 5117 11396 5173 11398
rect 4877 10362 4933 10364
rect 4957 10362 5013 10364
rect 5037 10362 5093 10364
rect 5117 10362 5173 10364
rect 4877 10310 4923 10362
rect 4923 10310 4933 10362
rect 4957 10310 4987 10362
rect 4987 10310 4999 10362
rect 4999 10310 5013 10362
rect 5037 10310 5051 10362
rect 5051 10310 5063 10362
rect 5063 10310 5093 10362
rect 5117 10310 5127 10362
rect 5127 10310 5173 10362
rect 4877 10308 4933 10310
rect 4957 10308 5013 10310
rect 5037 10308 5093 10310
rect 5117 10308 5173 10310
rect 4877 9274 4933 9276
rect 4957 9274 5013 9276
rect 5037 9274 5093 9276
rect 5117 9274 5173 9276
rect 4877 9222 4923 9274
rect 4923 9222 4933 9274
rect 4957 9222 4987 9274
rect 4987 9222 4999 9274
rect 4999 9222 5013 9274
rect 5037 9222 5051 9274
rect 5051 9222 5063 9274
rect 5063 9222 5093 9274
rect 5117 9222 5127 9274
rect 5127 9222 5173 9274
rect 4877 9220 4933 9222
rect 4957 9220 5013 9222
rect 5037 9220 5093 9222
rect 5117 9220 5173 9222
rect 5906 8880 5962 8936
rect 4877 8186 4933 8188
rect 4957 8186 5013 8188
rect 5037 8186 5093 8188
rect 5117 8186 5173 8188
rect 4877 8134 4923 8186
rect 4923 8134 4933 8186
rect 4957 8134 4987 8186
rect 4987 8134 4999 8186
rect 4999 8134 5013 8186
rect 5037 8134 5051 8186
rect 5051 8134 5063 8186
rect 5063 8134 5093 8186
rect 5117 8134 5127 8186
rect 5127 8134 5173 8186
rect 4877 8132 4933 8134
rect 4957 8132 5013 8134
rect 5037 8132 5093 8134
rect 5117 8132 5173 8134
rect 4877 7098 4933 7100
rect 4957 7098 5013 7100
rect 5037 7098 5093 7100
rect 5117 7098 5173 7100
rect 4877 7046 4923 7098
rect 4923 7046 4933 7098
rect 4957 7046 4987 7098
rect 4987 7046 4999 7098
rect 4999 7046 5013 7098
rect 5037 7046 5051 7098
rect 5051 7046 5063 7098
rect 5063 7046 5093 7098
rect 5117 7046 5127 7098
rect 5127 7046 5173 7098
rect 4877 7044 4933 7046
rect 4957 7044 5013 7046
rect 5037 7044 5093 7046
rect 5117 7044 5173 7046
rect 7746 17604 7802 17640
rect 7746 17584 7748 17604
rect 7748 17584 7800 17604
rect 7800 17584 7802 17604
rect 8798 18522 8854 18524
rect 8878 18522 8934 18524
rect 8958 18522 9014 18524
rect 9038 18522 9094 18524
rect 8798 18470 8844 18522
rect 8844 18470 8854 18522
rect 8878 18470 8908 18522
rect 8908 18470 8920 18522
rect 8920 18470 8934 18522
rect 8958 18470 8972 18522
rect 8972 18470 8984 18522
rect 8984 18470 9014 18522
rect 9038 18470 9048 18522
rect 9048 18470 9094 18522
rect 8798 18468 8854 18470
rect 8878 18468 8934 18470
rect 8958 18468 9014 18470
rect 9038 18468 9094 18470
rect 8798 17434 8854 17436
rect 8878 17434 8934 17436
rect 8958 17434 9014 17436
rect 9038 17434 9094 17436
rect 8798 17382 8844 17434
rect 8844 17382 8854 17434
rect 8878 17382 8908 17434
rect 8908 17382 8920 17434
rect 8920 17382 8934 17434
rect 8958 17382 8972 17434
rect 8972 17382 8984 17434
rect 8984 17382 9014 17434
rect 9038 17382 9048 17434
rect 9048 17382 9094 17434
rect 8798 17380 8854 17382
rect 8878 17380 8934 17382
rect 8958 17380 9014 17382
rect 9038 17380 9094 17382
rect 8798 16346 8854 16348
rect 8878 16346 8934 16348
rect 8958 16346 9014 16348
rect 9038 16346 9094 16348
rect 8798 16294 8844 16346
rect 8844 16294 8854 16346
rect 8878 16294 8908 16346
rect 8908 16294 8920 16346
rect 8920 16294 8934 16346
rect 8958 16294 8972 16346
rect 8972 16294 8984 16346
rect 8984 16294 9014 16346
rect 9038 16294 9048 16346
rect 9048 16294 9094 16346
rect 8798 16292 8854 16294
rect 8878 16292 8934 16294
rect 8958 16292 9014 16294
rect 9038 16292 9094 16294
rect 8798 15258 8854 15260
rect 8878 15258 8934 15260
rect 8958 15258 9014 15260
rect 9038 15258 9094 15260
rect 8798 15206 8844 15258
rect 8844 15206 8854 15258
rect 8878 15206 8908 15258
rect 8908 15206 8920 15258
rect 8920 15206 8934 15258
rect 8958 15206 8972 15258
rect 8972 15206 8984 15258
rect 8984 15206 9014 15258
rect 9038 15206 9048 15258
rect 9048 15206 9094 15258
rect 8798 15204 8854 15206
rect 8878 15204 8934 15206
rect 8958 15204 9014 15206
rect 9038 15204 9094 15206
rect 8666 14864 8722 14920
rect 8798 14170 8854 14172
rect 8878 14170 8934 14172
rect 8958 14170 9014 14172
rect 9038 14170 9094 14172
rect 8798 14118 8844 14170
rect 8844 14118 8854 14170
rect 8878 14118 8908 14170
rect 8908 14118 8920 14170
rect 8920 14118 8934 14170
rect 8958 14118 8972 14170
rect 8972 14118 8984 14170
rect 8984 14118 9014 14170
rect 9038 14118 9048 14170
rect 9048 14118 9094 14170
rect 8798 14116 8854 14118
rect 8878 14116 8934 14118
rect 8958 14116 9014 14118
rect 9038 14116 9094 14118
rect 8798 13082 8854 13084
rect 8878 13082 8934 13084
rect 8958 13082 9014 13084
rect 9038 13082 9094 13084
rect 8798 13030 8844 13082
rect 8844 13030 8854 13082
rect 8878 13030 8908 13082
rect 8908 13030 8920 13082
rect 8920 13030 8934 13082
rect 8958 13030 8972 13082
rect 8972 13030 8984 13082
rect 8984 13030 9014 13082
rect 9038 13030 9048 13082
rect 9048 13030 9094 13082
rect 8798 13028 8854 13030
rect 8878 13028 8934 13030
rect 8958 13028 9014 13030
rect 9038 13028 9094 13030
rect 9218 15952 9274 16008
rect 8798 11994 8854 11996
rect 8878 11994 8934 11996
rect 8958 11994 9014 11996
rect 9038 11994 9094 11996
rect 8798 11942 8844 11994
rect 8844 11942 8854 11994
rect 8878 11942 8908 11994
rect 8908 11942 8920 11994
rect 8920 11942 8934 11994
rect 8958 11942 8972 11994
rect 8972 11942 8984 11994
rect 8984 11942 9014 11994
rect 9038 11942 9048 11994
rect 9048 11942 9094 11994
rect 8798 11940 8854 11942
rect 8878 11940 8934 11942
rect 8958 11940 9014 11942
rect 9038 11940 9094 11942
rect 8798 10906 8854 10908
rect 8878 10906 8934 10908
rect 8958 10906 9014 10908
rect 9038 10906 9094 10908
rect 8798 10854 8844 10906
rect 8844 10854 8854 10906
rect 8878 10854 8908 10906
rect 8908 10854 8920 10906
rect 8920 10854 8934 10906
rect 8958 10854 8972 10906
rect 8972 10854 8984 10906
rect 8984 10854 9014 10906
rect 9038 10854 9048 10906
rect 9048 10854 9094 10906
rect 8798 10852 8854 10854
rect 8878 10852 8934 10854
rect 8958 10852 9014 10854
rect 9038 10852 9094 10854
rect 8798 9818 8854 9820
rect 8878 9818 8934 9820
rect 8958 9818 9014 9820
rect 9038 9818 9094 9820
rect 8798 9766 8844 9818
rect 8844 9766 8854 9818
rect 8878 9766 8908 9818
rect 8908 9766 8920 9818
rect 8920 9766 8934 9818
rect 8958 9766 8972 9818
rect 8972 9766 8984 9818
rect 8984 9766 9014 9818
rect 9038 9766 9048 9818
rect 9048 9766 9094 9818
rect 8798 9764 8854 9766
rect 8878 9764 8934 9766
rect 8958 9764 9014 9766
rect 9038 9764 9094 9766
rect 8798 8730 8854 8732
rect 8878 8730 8934 8732
rect 8958 8730 9014 8732
rect 9038 8730 9094 8732
rect 8798 8678 8844 8730
rect 8844 8678 8854 8730
rect 8878 8678 8908 8730
rect 8908 8678 8920 8730
rect 8920 8678 8934 8730
rect 8958 8678 8972 8730
rect 8972 8678 8984 8730
rect 8984 8678 9014 8730
rect 9038 8678 9048 8730
rect 9048 8678 9094 8730
rect 8798 8676 8854 8678
rect 8878 8676 8934 8678
rect 8958 8676 9014 8678
rect 9038 8676 9094 8678
rect 8798 7642 8854 7644
rect 8878 7642 8934 7644
rect 8958 7642 9014 7644
rect 9038 7642 9094 7644
rect 8798 7590 8844 7642
rect 8844 7590 8854 7642
rect 8878 7590 8908 7642
rect 8908 7590 8920 7642
rect 8920 7590 8934 7642
rect 8958 7590 8972 7642
rect 8972 7590 8984 7642
rect 8984 7590 9014 7642
rect 9038 7590 9048 7642
rect 9048 7590 9094 7642
rect 8798 7588 8854 7590
rect 8878 7588 8934 7590
rect 8958 7588 9014 7590
rect 9038 7588 9094 7590
rect 9586 16124 9588 16144
rect 9588 16124 9640 16144
rect 9640 16124 9642 16144
rect 9586 16088 9642 16124
rect 10414 16652 10470 16688
rect 10414 16632 10416 16652
rect 10416 16632 10468 16652
rect 10468 16632 10470 16652
rect 11150 18692 11206 18728
rect 11150 18672 11152 18692
rect 11152 18672 11204 18692
rect 11204 18672 11206 18692
rect 13082 21120 13138 21176
rect 11058 17196 11114 17232
rect 11058 17176 11060 17196
rect 11060 17176 11112 17196
rect 11112 17176 11114 17196
rect 11702 17756 11704 17776
rect 11704 17756 11756 17776
rect 11756 17756 11758 17776
rect 11702 17720 11758 17756
rect 12719 20154 12775 20156
rect 12799 20154 12855 20156
rect 12879 20154 12935 20156
rect 12959 20154 13015 20156
rect 12719 20102 12765 20154
rect 12765 20102 12775 20154
rect 12799 20102 12829 20154
rect 12829 20102 12841 20154
rect 12841 20102 12855 20154
rect 12879 20102 12893 20154
rect 12893 20102 12905 20154
rect 12905 20102 12935 20154
rect 12959 20102 12969 20154
rect 12969 20102 13015 20154
rect 12719 20100 12775 20102
rect 12799 20100 12855 20102
rect 12879 20100 12935 20102
rect 12959 20100 13015 20102
rect 12346 18128 12402 18184
rect 13542 20596 13598 20632
rect 13542 20576 13544 20596
rect 13544 20576 13596 20596
rect 13596 20576 13598 20596
rect 12719 19066 12775 19068
rect 12799 19066 12855 19068
rect 12879 19066 12935 19068
rect 12959 19066 13015 19068
rect 12719 19014 12765 19066
rect 12765 19014 12775 19066
rect 12799 19014 12829 19066
rect 12829 19014 12841 19066
rect 12841 19014 12855 19066
rect 12879 19014 12893 19066
rect 12893 19014 12905 19066
rect 12905 19014 12935 19066
rect 12959 19014 12969 19066
rect 12969 19014 13015 19066
rect 12719 19012 12775 19014
rect 12799 19012 12855 19014
rect 12879 19012 12935 19014
rect 12959 19012 13015 19014
rect 12719 17978 12775 17980
rect 12799 17978 12855 17980
rect 12879 17978 12935 17980
rect 12959 17978 13015 17980
rect 12719 17926 12765 17978
rect 12765 17926 12775 17978
rect 12799 17926 12829 17978
rect 12829 17926 12841 17978
rect 12841 17926 12855 17978
rect 12879 17926 12893 17978
rect 12893 17926 12905 17978
rect 12905 17926 12935 17978
rect 12959 17926 12969 17978
rect 12969 17926 13015 17978
rect 12719 17924 12775 17926
rect 12799 17924 12855 17926
rect 12879 17924 12935 17926
rect 12959 17924 13015 17926
rect 11518 13368 11574 13424
rect 9678 9580 9734 9616
rect 9678 9560 9680 9580
rect 9680 9560 9732 9580
rect 9732 9560 9734 9580
rect 8798 6554 8854 6556
rect 8878 6554 8934 6556
rect 8958 6554 9014 6556
rect 9038 6554 9094 6556
rect 8798 6502 8844 6554
rect 8844 6502 8854 6554
rect 8878 6502 8908 6554
rect 8908 6502 8920 6554
rect 8920 6502 8934 6554
rect 8958 6502 8972 6554
rect 8972 6502 8984 6554
rect 8984 6502 9014 6554
rect 9038 6502 9048 6554
rect 9048 6502 9094 6554
rect 8798 6500 8854 6502
rect 8878 6500 8934 6502
rect 8958 6500 9014 6502
rect 9038 6500 9094 6502
rect 10414 9580 10470 9616
rect 10414 9560 10416 9580
rect 10416 9560 10468 9580
rect 10468 9560 10470 9580
rect 10138 8472 10194 8528
rect 13358 18708 13360 18728
rect 13360 18708 13412 18728
rect 13412 18708 13414 18728
rect 13358 18672 13414 18708
rect 13082 17448 13138 17504
rect 12719 16890 12775 16892
rect 12799 16890 12855 16892
rect 12879 16890 12935 16892
rect 12959 16890 13015 16892
rect 12719 16838 12765 16890
rect 12765 16838 12775 16890
rect 12799 16838 12829 16890
rect 12829 16838 12841 16890
rect 12841 16838 12855 16890
rect 12879 16838 12893 16890
rect 12893 16838 12905 16890
rect 12905 16838 12935 16890
rect 12959 16838 12969 16890
rect 12969 16838 13015 16890
rect 12719 16836 12775 16838
rect 12799 16836 12855 16838
rect 12879 16836 12935 16838
rect 12959 16836 13015 16838
rect 27342 20984 27398 21040
rect 17130 20848 17186 20904
rect 16640 20698 16696 20700
rect 16720 20698 16776 20700
rect 16800 20698 16856 20700
rect 16880 20698 16936 20700
rect 16640 20646 16686 20698
rect 16686 20646 16696 20698
rect 16720 20646 16750 20698
rect 16750 20646 16762 20698
rect 16762 20646 16776 20698
rect 16800 20646 16814 20698
rect 16814 20646 16826 20698
rect 16826 20646 16856 20698
rect 16880 20646 16890 20698
rect 16890 20646 16936 20698
rect 16640 20644 16696 20646
rect 16720 20644 16776 20646
rect 16800 20644 16856 20646
rect 16880 20644 16936 20646
rect 16118 20596 16174 20632
rect 16118 20576 16120 20596
rect 16120 20576 16172 20596
rect 16172 20576 16174 20596
rect 17038 20596 17094 20632
rect 17038 20576 17040 20596
rect 17040 20576 17092 20596
rect 17092 20576 17094 20596
rect 13726 19352 13782 19408
rect 14186 18128 14242 18184
rect 13082 16108 13138 16144
rect 13082 16088 13084 16108
rect 13084 16088 13136 16108
rect 13136 16088 13138 16108
rect 12719 15802 12775 15804
rect 12799 15802 12855 15804
rect 12879 15802 12935 15804
rect 12959 15802 13015 15804
rect 12719 15750 12765 15802
rect 12765 15750 12775 15802
rect 12799 15750 12829 15802
rect 12829 15750 12841 15802
rect 12841 15750 12855 15802
rect 12879 15750 12893 15802
rect 12893 15750 12905 15802
rect 12905 15750 12935 15802
rect 12959 15750 12969 15802
rect 12969 15750 13015 15802
rect 12719 15748 12775 15750
rect 12799 15748 12855 15750
rect 12879 15748 12935 15750
rect 12959 15748 13015 15750
rect 12719 14714 12775 14716
rect 12799 14714 12855 14716
rect 12879 14714 12935 14716
rect 12959 14714 13015 14716
rect 12719 14662 12765 14714
rect 12765 14662 12775 14714
rect 12799 14662 12829 14714
rect 12829 14662 12841 14714
rect 12841 14662 12855 14714
rect 12879 14662 12893 14714
rect 12893 14662 12905 14714
rect 12905 14662 12935 14714
rect 12959 14662 12969 14714
rect 12969 14662 13015 14714
rect 12719 14660 12775 14662
rect 12799 14660 12855 14662
rect 12879 14660 12935 14662
rect 12959 14660 13015 14662
rect 12714 14456 12770 14512
rect 13082 13912 13138 13968
rect 12719 13626 12775 13628
rect 12799 13626 12855 13628
rect 12879 13626 12935 13628
rect 12959 13626 13015 13628
rect 12719 13574 12765 13626
rect 12765 13574 12775 13626
rect 12799 13574 12829 13626
rect 12829 13574 12841 13626
rect 12841 13574 12855 13626
rect 12879 13574 12893 13626
rect 12893 13574 12905 13626
rect 12905 13574 12935 13626
rect 12959 13574 12969 13626
rect 12969 13574 13015 13626
rect 12719 13572 12775 13574
rect 12799 13572 12855 13574
rect 12879 13572 12935 13574
rect 12959 13572 13015 13574
rect 12719 12538 12775 12540
rect 12799 12538 12855 12540
rect 12879 12538 12935 12540
rect 12959 12538 13015 12540
rect 12719 12486 12765 12538
rect 12765 12486 12775 12538
rect 12799 12486 12829 12538
rect 12829 12486 12841 12538
rect 12841 12486 12855 12538
rect 12879 12486 12893 12538
rect 12893 12486 12905 12538
rect 12905 12486 12935 12538
rect 12959 12486 12969 12538
rect 12969 12486 13015 12538
rect 12719 12484 12775 12486
rect 12799 12484 12855 12486
rect 12879 12484 12935 12486
rect 12959 12484 13015 12486
rect 11426 9560 11482 9616
rect 12719 11450 12775 11452
rect 12799 11450 12855 11452
rect 12879 11450 12935 11452
rect 12959 11450 13015 11452
rect 12719 11398 12765 11450
rect 12765 11398 12775 11450
rect 12799 11398 12829 11450
rect 12829 11398 12841 11450
rect 12841 11398 12855 11450
rect 12879 11398 12893 11450
rect 12893 11398 12905 11450
rect 12905 11398 12935 11450
rect 12959 11398 12969 11450
rect 12969 11398 13015 11450
rect 12719 11396 12775 11398
rect 12799 11396 12855 11398
rect 12879 11396 12935 11398
rect 12959 11396 13015 11398
rect 13726 15000 13782 15056
rect 14554 17720 14610 17776
rect 14830 16532 14832 16552
rect 14832 16532 14884 16552
rect 14884 16532 14886 16552
rect 14830 16496 14886 16532
rect 14370 14456 14426 14512
rect 13174 12960 13230 13016
rect 12719 10362 12775 10364
rect 12799 10362 12855 10364
rect 12879 10362 12935 10364
rect 12959 10362 13015 10364
rect 12719 10310 12765 10362
rect 12765 10310 12775 10362
rect 12799 10310 12829 10362
rect 12829 10310 12841 10362
rect 12841 10310 12855 10362
rect 12879 10310 12893 10362
rect 12893 10310 12905 10362
rect 12905 10310 12935 10362
rect 12959 10310 12969 10362
rect 12969 10310 13015 10362
rect 12719 10308 12775 10310
rect 12799 10308 12855 10310
rect 12879 10308 12935 10310
rect 12959 10308 13015 10310
rect 12719 9274 12775 9276
rect 12799 9274 12855 9276
rect 12879 9274 12935 9276
rect 12959 9274 13015 9276
rect 12719 9222 12765 9274
rect 12765 9222 12775 9274
rect 12799 9222 12829 9274
rect 12829 9222 12841 9274
rect 12841 9222 12855 9274
rect 12879 9222 12893 9274
rect 12893 9222 12905 9274
rect 12905 9222 12935 9274
rect 12959 9222 12969 9274
rect 12969 9222 13015 9274
rect 12719 9220 12775 9222
rect 12799 9220 12855 9222
rect 12879 9220 12935 9222
rect 12959 9220 13015 9222
rect 14278 12316 14280 12336
rect 14280 12316 14332 12336
rect 14332 12316 14334 12336
rect 14278 12280 14334 12316
rect 14646 13232 14702 13288
rect 14738 12960 14794 13016
rect 14462 11756 14518 11792
rect 14462 11736 14464 11756
rect 14464 11736 14516 11756
rect 14516 11736 14518 11756
rect 13634 11056 13690 11112
rect 13542 9560 13598 9616
rect 12719 8186 12775 8188
rect 12799 8186 12855 8188
rect 12879 8186 12935 8188
rect 12959 8186 13015 8188
rect 12719 8134 12765 8186
rect 12765 8134 12775 8186
rect 12799 8134 12829 8186
rect 12829 8134 12841 8186
rect 12841 8134 12855 8186
rect 12879 8134 12893 8186
rect 12893 8134 12905 8186
rect 12905 8134 12935 8186
rect 12959 8134 12969 8186
rect 12969 8134 13015 8186
rect 12719 8132 12775 8134
rect 12799 8132 12855 8134
rect 12879 8132 12935 8134
rect 12959 8132 13015 8134
rect 12719 7098 12775 7100
rect 12799 7098 12855 7100
rect 12879 7098 12935 7100
rect 12959 7098 13015 7100
rect 12719 7046 12765 7098
rect 12765 7046 12775 7098
rect 12799 7046 12829 7098
rect 12829 7046 12841 7098
rect 12841 7046 12855 7098
rect 12879 7046 12893 7098
rect 12893 7046 12905 7098
rect 12905 7046 12935 7098
rect 12959 7046 12969 7098
rect 12969 7046 13015 7098
rect 12719 7044 12775 7046
rect 12799 7044 12855 7046
rect 12879 7044 12935 7046
rect 12959 7044 13015 7046
rect 13634 8880 13690 8936
rect 15014 17856 15070 17912
rect 15106 17448 15162 17504
rect 15474 17856 15530 17912
rect 15198 16904 15254 16960
rect 16640 19610 16696 19612
rect 16720 19610 16776 19612
rect 16800 19610 16856 19612
rect 16880 19610 16936 19612
rect 16640 19558 16686 19610
rect 16686 19558 16696 19610
rect 16720 19558 16750 19610
rect 16750 19558 16762 19610
rect 16762 19558 16776 19610
rect 16800 19558 16814 19610
rect 16814 19558 16826 19610
rect 16826 19558 16856 19610
rect 16880 19558 16890 19610
rect 16890 19558 16936 19610
rect 16640 19556 16696 19558
rect 16720 19556 16776 19558
rect 16800 19556 16856 19558
rect 16880 19556 16936 19558
rect 24482 20698 24538 20700
rect 24562 20698 24618 20700
rect 24642 20698 24698 20700
rect 24722 20698 24778 20700
rect 24482 20646 24528 20698
rect 24528 20646 24538 20698
rect 24562 20646 24592 20698
rect 24592 20646 24604 20698
rect 24604 20646 24618 20698
rect 24642 20646 24656 20698
rect 24656 20646 24668 20698
rect 24668 20646 24698 20698
rect 24722 20646 24732 20698
rect 24732 20646 24778 20698
rect 24482 20644 24538 20646
rect 24562 20644 24618 20646
rect 24642 20644 24698 20646
rect 24722 20644 24778 20646
rect 16210 17856 16266 17912
rect 16640 18522 16696 18524
rect 16720 18522 16776 18524
rect 16800 18522 16856 18524
rect 16880 18522 16936 18524
rect 16640 18470 16686 18522
rect 16686 18470 16696 18522
rect 16720 18470 16750 18522
rect 16750 18470 16762 18522
rect 16762 18470 16776 18522
rect 16800 18470 16814 18522
rect 16814 18470 16826 18522
rect 16826 18470 16856 18522
rect 16880 18470 16890 18522
rect 16890 18470 16936 18522
rect 16640 18468 16696 18470
rect 16720 18468 16776 18470
rect 16800 18468 16856 18470
rect 16880 18468 16936 18470
rect 16640 17434 16696 17436
rect 16720 17434 16776 17436
rect 16800 17434 16856 17436
rect 16880 17434 16936 17436
rect 16640 17382 16686 17434
rect 16686 17382 16696 17434
rect 16720 17382 16750 17434
rect 16750 17382 16762 17434
rect 16762 17382 16776 17434
rect 16800 17382 16814 17434
rect 16814 17382 16826 17434
rect 16826 17382 16856 17434
rect 16880 17382 16890 17434
rect 16890 17382 16936 17434
rect 16640 17380 16696 17382
rect 16720 17380 16776 17382
rect 16800 17380 16856 17382
rect 16880 17380 16936 17382
rect 16394 16632 16450 16688
rect 14186 8492 14242 8528
rect 14186 8472 14188 8492
rect 14188 8472 14240 8492
rect 14240 8472 14242 8492
rect 4877 6010 4933 6012
rect 4957 6010 5013 6012
rect 5037 6010 5093 6012
rect 5117 6010 5173 6012
rect 4877 5958 4923 6010
rect 4923 5958 4933 6010
rect 4957 5958 4987 6010
rect 4987 5958 4999 6010
rect 4999 5958 5013 6010
rect 5037 5958 5051 6010
rect 5051 5958 5063 6010
rect 5063 5958 5093 6010
rect 5117 5958 5127 6010
rect 5127 5958 5173 6010
rect 4877 5956 4933 5958
rect 4957 5956 5013 5958
rect 5037 5956 5093 5958
rect 5117 5956 5173 5958
rect 12719 6010 12775 6012
rect 12799 6010 12855 6012
rect 12879 6010 12935 6012
rect 12959 6010 13015 6012
rect 12719 5958 12765 6010
rect 12765 5958 12775 6010
rect 12799 5958 12829 6010
rect 12829 5958 12841 6010
rect 12841 5958 12855 6010
rect 12879 5958 12893 6010
rect 12893 5958 12905 6010
rect 12905 5958 12935 6010
rect 12959 5958 12969 6010
rect 12969 5958 13015 6010
rect 12719 5956 12775 5958
rect 12799 5956 12855 5958
rect 12879 5956 12935 5958
rect 12959 5956 13015 5958
rect 15566 12960 15622 13016
rect 18602 19508 18658 19544
rect 18602 19488 18604 19508
rect 18604 19488 18656 19508
rect 18656 19488 18658 19508
rect 19614 19216 19670 19272
rect 17590 17040 17646 17096
rect 16640 16346 16696 16348
rect 16720 16346 16776 16348
rect 16800 16346 16856 16348
rect 16880 16346 16936 16348
rect 16640 16294 16686 16346
rect 16686 16294 16696 16346
rect 16720 16294 16750 16346
rect 16750 16294 16762 16346
rect 16762 16294 16776 16346
rect 16800 16294 16814 16346
rect 16814 16294 16826 16346
rect 16826 16294 16856 16346
rect 16880 16294 16890 16346
rect 16890 16294 16936 16346
rect 16640 16292 16696 16294
rect 16720 16292 16776 16294
rect 16800 16292 16856 16294
rect 16880 16292 16936 16294
rect 18510 16904 18566 16960
rect 18786 16904 18842 16960
rect 18418 16360 18474 16416
rect 16640 15258 16696 15260
rect 16720 15258 16776 15260
rect 16800 15258 16856 15260
rect 16880 15258 16936 15260
rect 16640 15206 16686 15258
rect 16686 15206 16696 15258
rect 16720 15206 16750 15258
rect 16750 15206 16762 15258
rect 16762 15206 16776 15258
rect 16800 15206 16814 15258
rect 16814 15206 16826 15258
rect 16826 15206 16856 15258
rect 16880 15206 16890 15258
rect 16890 15206 16936 15258
rect 16640 15204 16696 15206
rect 16720 15204 16776 15206
rect 16800 15204 16856 15206
rect 16880 15204 16936 15206
rect 16640 14170 16696 14172
rect 16720 14170 16776 14172
rect 16800 14170 16856 14172
rect 16880 14170 16936 14172
rect 16640 14118 16686 14170
rect 16686 14118 16696 14170
rect 16720 14118 16750 14170
rect 16750 14118 16762 14170
rect 16762 14118 16776 14170
rect 16800 14118 16814 14170
rect 16814 14118 16826 14170
rect 16826 14118 16856 14170
rect 16880 14118 16890 14170
rect 16890 14118 16936 14170
rect 16640 14116 16696 14118
rect 16720 14116 16776 14118
rect 16800 14116 16856 14118
rect 16880 14116 16936 14118
rect 16640 13082 16696 13084
rect 16720 13082 16776 13084
rect 16800 13082 16856 13084
rect 16880 13082 16936 13084
rect 16640 13030 16686 13082
rect 16686 13030 16696 13082
rect 16720 13030 16750 13082
rect 16750 13030 16762 13082
rect 16762 13030 16776 13082
rect 16800 13030 16814 13082
rect 16814 13030 16826 13082
rect 16826 13030 16856 13082
rect 16880 13030 16890 13082
rect 16890 13030 16936 13082
rect 16640 13028 16696 13030
rect 16720 13028 16776 13030
rect 16800 13028 16856 13030
rect 16880 13028 16936 13030
rect 20561 20154 20617 20156
rect 20641 20154 20697 20156
rect 20721 20154 20777 20156
rect 20801 20154 20857 20156
rect 20561 20102 20607 20154
rect 20607 20102 20617 20154
rect 20641 20102 20671 20154
rect 20671 20102 20683 20154
rect 20683 20102 20697 20154
rect 20721 20102 20735 20154
rect 20735 20102 20747 20154
rect 20747 20102 20777 20154
rect 20801 20102 20811 20154
rect 20811 20102 20857 20154
rect 20561 20100 20617 20102
rect 20641 20100 20697 20102
rect 20721 20100 20777 20102
rect 20801 20100 20857 20102
rect 20561 19066 20617 19068
rect 20641 19066 20697 19068
rect 20721 19066 20777 19068
rect 20801 19066 20857 19068
rect 20561 19014 20607 19066
rect 20607 19014 20617 19066
rect 20641 19014 20671 19066
rect 20671 19014 20683 19066
rect 20683 19014 20697 19066
rect 20721 19014 20735 19066
rect 20735 19014 20747 19066
rect 20747 19014 20777 19066
rect 20801 19014 20811 19066
rect 20811 19014 20857 19066
rect 20561 19012 20617 19014
rect 20641 19012 20697 19014
rect 20721 19012 20777 19014
rect 20801 19012 20857 19014
rect 20561 17978 20617 17980
rect 20641 17978 20697 17980
rect 20721 17978 20777 17980
rect 20801 17978 20857 17980
rect 20561 17926 20607 17978
rect 20607 17926 20617 17978
rect 20641 17926 20671 17978
rect 20671 17926 20683 17978
rect 20683 17926 20697 17978
rect 20721 17926 20735 17978
rect 20735 17926 20747 17978
rect 20747 17926 20777 17978
rect 20801 17926 20811 17978
rect 20811 17926 20857 17978
rect 20561 17924 20617 17926
rect 20641 17924 20697 17926
rect 20721 17924 20777 17926
rect 20801 17924 20857 17926
rect 19246 16496 19302 16552
rect 20561 16890 20617 16892
rect 20641 16890 20697 16892
rect 20721 16890 20777 16892
rect 20801 16890 20857 16892
rect 20561 16838 20607 16890
rect 20607 16838 20617 16890
rect 20641 16838 20671 16890
rect 20671 16838 20683 16890
rect 20683 16838 20697 16890
rect 20721 16838 20735 16890
rect 20735 16838 20747 16890
rect 20747 16838 20777 16890
rect 20801 16838 20811 16890
rect 20811 16838 20857 16890
rect 20561 16836 20617 16838
rect 20641 16836 20697 16838
rect 20721 16836 20777 16838
rect 20801 16836 20857 16838
rect 21086 17856 21142 17912
rect 20994 17176 21050 17232
rect 21178 16516 21234 16552
rect 21178 16496 21180 16516
rect 21180 16496 21232 16516
rect 21232 16496 21234 16516
rect 19982 16088 20038 16144
rect 20994 16360 21050 16416
rect 20561 15802 20617 15804
rect 20641 15802 20697 15804
rect 20721 15802 20777 15804
rect 20801 15802 20857 15804
rect 20561 15750 20607 15802
rect 20607 15750 20617 15802
rect 20641 15750 20671 15802
rect 20671 15750 20683 15802
rect 20683 15750 20697 15802
rect 20721 15750 20735 15802
rect 20735 15750 20747 15802
rect 20747 15750 20777 15802
rect 20801 15750 20811 15802
rect 20811 15750 20857 15802
rect 20561 15748 20617 15750
rect 20641 15748 20697 15750
rect 20721 15748 20777 15750
rect 20801 15748 20857 15750
rect 19982 15408 20038 15464
rect 18418 13912 18474 13968
rect 16640 11994 16696 11996
rect 16720 11994 16776 11996
rect 16800 11994 16856 11996
rect 16880 11994 16936 11996
rect 16640 11942 16686 11994
rect 16686 11942 16696 11994
rect 16720 11942 16750 11994
rect 16750 11942 16762 11994
rect 16762 11942 16776 11994
rect 16800 11942 16814 11994
rect 16814 11942 16826 11994
rect 16826 11942 16856 11994
rect 16880 11942 16890 11994
rect 16890 11942 16936 11994
rect 16640 11940 16696 11942
rect 16720 11940 16776 11942
rect 16800 11940 16856 11942
rect 16880 11940 16936 11942
rect 20561 14714 20617 14716
rect 20641 14714 20697 14716
rect 20721 14714 20777 14716
rect 20801 14714 20857 14716
rect 20561 14662 20607 14714
rect 20607 14662 20617 14714
rect 20641 14662 20671 14714
rect 20671 14662 20683 14714
rect 20683 14662 20697 14714
rect 20721 14662 20735 14714
rect 20735 14662 20747 14714
rect 20747 14662 20777 14714
rect 20801 14662 20811 14714
rect 20811 14662 20857 14714
rect 20561 14660 20617 14662
rect 20641 14660 20697 14662
rect 20721 14660 20777 14662
rect 20801 14660 20857 14662
rect 20166 13776 20222 13832
rect 20561 13626 20617 13628
rect 20641 13626 20697 13628
rect 20721 13626 20777 13628
rect 20801 13626 20857 13628
rect 20561 13574 20607 13626
rect 20607 13574 20617 13626
rect 20641 13574 20671 13626
rect 20671 13574 20683 13626
rect 20683 13574 20697 13626
rect 20721 13574 20735 13626
rect 20735 13574 20747 13626
rect 20747 13574 20777 13626
rect 20801 13574 20811 13626
rect 20811 13574 20857 13626
rect 20561 13572 20617 13574
rect 20641 13572 20697 13574
rect 20721 13572 20777 13574
rect 20801 13572 20857 13574
rect 21270 15136 21326 15192
rect 21638 15444 21640 15464
rect 21640 15444 21692 15464
rect 21692 15444 21694 15464
rect 21638 15408 21694 15444
rect 21914 15272 21970 15328
rect 20561 12538 20617 12540
rect 20641 12538 20697 12540
rect 20721 12538 20777 12540
rect 20801 12538 20857 12540
rect 20561 12486 20607 12538
rect 20607 12486 20617 12538
rect 20641 12486 20671 12538
rect 20671 12486 20683 12538
rect 20683 12486 20697 12538
rect 20721 12486 20735 12538
rect 20735 12486 20747 12538
rect 20747 12486 20777 12538
rect 20801 12486 20811 12538
rect 20811 12486 20857 12538
rect 20561 12484 20617 12486
rect 20641 12484 20697 12486
rect 20721 12484 20777 12486
rect 20801 12484 20857 12486
rect 16946 11076 17002 11112
rect 16946 11056 16948 11076
rect 16948 11056 17000 11076
rect 17000 11056 17002 11076
rect 16640 10906 16696 10908
rect 16720 10906 16776 10908
rect 16800 10906 16856 10908
rect 16880 10906 16936 10908
rect 16640 10854 16686 10906
rect 16686 10854 16696 10906
rect 16720 10854 16750 10906
rect 16750 10854 16762 10906
rect 16762 10854 16776 10906
rect 16800 10854 16814 10906
rect 16814 10854 16826 10906
rect 16826 10854 16856 10906
rect 16880 10854 16890 10906
rect 16890 10854 16936 10906
rect 16640 10852 16696 10854
rect 16720 10852 16776 10854
rect 16800 10852 16856 10854
rect 16880 10852 16936 10854
rect 16640 9818 16696 9820
rect 16720 9818 16776 9820
rect 16800 9818 16856 9820
rect 16880 9818 16936 9820
rect 16640 9766 16686 9818
rect 16686 9766 16696 9818
rect 16720 9766 16750 9818
rect 16750 9766 16762 9818
rect 16762 9766 16776 9818
rect 16800 9766 16814 9818
rect 16814 9766 16826 9818
rect 16826 9766 16856 9818
rect 16880 9766 16890 9818
rect 16890 9766 16936 9818
rect 16640 9764 16696 9766
rect 16720 9764 16776 9766
rect 16800 9764 16856 9766
rect 16880 9764 16936 9766
rect 18786 11756 18842 11792
rect 18786 11736 18788 11756
rect 18788 11736 18840 11756
rect 18840 11736 18842 11756
rect 20561 11450 20617 11452
rect 20641 11450 20697 11452
rect 20721 11450 20777 11452
rect 20801 11450 20857 11452
rect 20561 11398 20607 11450
rect 20607 11398 20617 11450
rect 20641 11398 20671 11450
rect 20671 11398 20683 11450
rect 20683 11398 20697 11450
rect 20721 11398 20735 11450
rect 20735 11398 20747 11450
rect 20747 11398 20777 11450
rect 20801 11398 20811 11450
rect 20811 11398 20857 11450
rect 20561 11396 20617 11398
rect 20641 11396 20697 11398
rect 20721 11396 20777 11398
rect 20801 11396 20857 11398
rect 16640 8730 16696 8732
rect 16720 8730 16776 8732
rect 16800 8730 16856 8732
rect 16880 8730 16936 8732
rect 16640 8678 16686 8730
rect 16686 8678 16696 8730
rect 16720 8678 16750 8730
rect 16750 8678 16762 8730
rect 16762 8678 16776 8730
rect 16800 8678 16814 8730
rect 16814 8678 16826 8730
rect 16826 8678 16856 8730
rect 16880 8678 16890 8730
rect 16890 8678 16936 8730
rect 16640 8676 16696 8678
rect 16720 8676 16776 8678
rect 16800 8676 16856 8678
rect 16880 8676 16936 8678
rect 16640 7642 16696 7644
rect 16720 7642 16776 7644
rect 16800 7642 16856 7644
rect 16880 7642 16936 7644
rect 16640 7590 16686 7642
rect 16686 7590 16696 7642
rect 16720 7590 16750 7642
rect 16750 7590 16762 7642
rect 16762 7590 16776 7642
rect 16800 7590 16814 7642
rect 16814 7590 16826 7642
rect 16826 7590 16856 7642
rect 16880 7590 16890 7642
rect 16890 7590 16936 7642
rect 16640 7588 16696 7590
rect 16720 7588 16776 7590
rect 16800 7588 16856 7590
rect 16880 7588 16936 7590
rect 16640 6554 16696 6556
rect 16720 6554 16776 6556
rect 16800 6554 16856 6556
rect 16880 6554 16936 6556
rect 16640 6502 16686 6554
rect 16686 6502 16696 6554
rect 16720 6502 16750 6554
rect 16750 6502 16762 6554
rect 16762 6502 16776 6554
rect 16800 6502 16814 6554
rect 16814 6502 16826 6554
rect 16826 6502 16856 6554
rect 16880 6502 16890 6554
rect 16890 6502 16936 6554
rect 16640 6500 16696 6502
rect 16720 6500 16776 6502
rect 16800 6500 16856 6502
rect 16880 6500 16936 6502
rect 8798 5466 8854 5468
rect 8878 5466 8934 5468
rect 8958 5466 9014 5468
rect 9038 5466 9094 5468
rect 8798 5414 8844 5466
rect 8844 5414 8854 5466
rect 8878 5414 8908 5466
rect 8908 5414 8920 5466
rect 8920 5414 8934 5466
rect 8958 5414 8972 5466
rect 8972 5414 8984 5466
rect 8984 5414 9014 5466
rect 9038 5414 9048 5466
rect 9048 5414 9094 5466
rect 8798 5412 8854 5414
rect 8878 5412 8934 5414
rect 8958 5412 9014 5414
rect 9038 5412 9094 5414
rect 16640 5466 16696 5468
rect 16720 5466 16776 5468
rect 16800 5466 16856 5468
rect 16880 5466 16936 5468
rect 16640 5414 16686 5466
rect 16686 5414 16696 5466
rect 16720 5414 16750 5466
rect 16750 5414 16762 5466
rect 16762 5414 16776 5466
rect 16800 5414 16814 5466
rect 16814 5414 16826 5466
rect 16826 5414 16856 5466
rect 16880 5414 16890 5466
rect 16890 5414 16936 5466
rect 16640 5412 16696 5414
rect 16720 5412 16776 5414
rect 16800 5412 16856 5414
rect 16880 5412 16936 5414
rect 20561 10362 20617 10364
rect 20641 10362 20697 10364
rect 20721 10362 20777 10364
rect 20801 10362 20857 10364
rect 20561 10310 20607 10362
rect 20607 10310 20617 10362
rect 20641 10310 20671 10362
rect 20671 10310 20683 10362
rect 20683 10310 20697 10362
rect 20721 10310 20735 10362
rect 20735 10310 20747 10362
rect 20747 10310 20777 10362
rect 20801 10310 20811 10362
rect 20811 10310 20857 10362
rect 20561 10308 20617 10310
rect 20641 10308 20697 10310
rect 20721 10308 20777 10310
rect 20801 10308 20857 10310
rect 22282 19252 22284 19272
rect 22284 19252 22336 19272
rect 22336 19252 22338 19272
rect 22282 19216 22338 19252
rect 24482 19610 24538 19612
rect 24562 19610 24618 19612
rect 24642 19610 24698 19612
rect 24722 19610 24778 19612
rect 24482 19558 24528 19610
rect 24528 19558 24538 19610
rect 24562 19558 24592 19610
rect 24592 19558 24604 19610
rect 24604 19558 24618 19610
rect 24642 19558 24656 19610
rect 24656 19558 24668 19610
rect 24668 19558 24698 19610
rect 24722 19558 24732 19610
rect 24732 19558 24778 19610
rect 24482 19556 24538 19558
rect 24562 19556 24618 19558
rect 24642 19556 24698 19558
rect 24722 19556 24778 19558
rect 24482 18522 24538 18524
rect 24562 18522 24618 18524
rect 24642 18522 24698 18524
rect 24722 18522 24778 18524
rect 24482 18470 24528 18522
rect 24528 18470 24538 18522
rect 24562 18470 24592 18522
rect 24592 18470 24604 18522
rect 24604 18470 24618 18522
rect 24642 18470 24656 18522
rect 24656 18470 24668 18522
rect 24668 18470 24698 18522
rect 24722 18470 24732 18522
rect 24732 18470 24778 18522
rect 24482 18468 24538 18470
rect 24562 18468 24618 18470
rect 24642 18468 24698 18470
rect 24722 18468 24778 18470
rect 22190 14864 22246 14920
rect 22006 13368 22062 13424
rect 23478 15444 23480 15464
rect 23480 15444 23532 15464
rect 23532 15444 23534 15464
rect 23478 15408 23534 15444
rect 23662 16496 23718 16552
rect 23754 16088 23810 16144
rect 23662 15272 23718 15328
rect 23662 15136 23718 15192
rect 20561 9274 20617 9276
rect 20641 9274 20697 9276
rect 20721 9274 20777 9276
rect 20801 9274 20857 9276
rect 20561 9222 20607 9274
rect 20607 9222 20617 9274
rect 20641 9222 20671 9274
rect 20671 9222 20683 9274
rect 20683 9222 20697 9274
rect 20721 9222 20735 9274
rect 20735 9222 20747 9274
rect 20747 9222 20777 9274
rect 20801 9222 20811 9274
rect 20811 9222 20857 9274
rect 20561 9220 20617 9222
rect 20641 9220 20697 9222
rect 20721 9220 20777 9222
rect 20801 9220 20857 9222
rect 20718 9016 20774 9072
rect 20561 8186 20617 8188
rect 20641 8186 20697 8188
rect 20721 8186 20777 8188
rect 20801 8186 20857 8188
rect 20561 8134 20607 8186
rect 20607 8134 20617 8186
rect 20641 8134 20671 8186
rect 20671 8134 20683 8186
rect 20683 8134 20697 8186
rect 20721 8134 20735 8186
rect 20735 8134 20747 8186
rect 20747 8134 20777 8186
rect 20801 8134 20811 8186
rect 20811 8134 20857 8186
rect 20561 8132 20617 8134
rect 20641 8132 20697 8134
rect 20721 8132 20777 8134
rect 20801 8132 20857 8134
rect 20561 7098 20617 7100
rect 20641 7098 20697 7100
rect 20721 7098 20777 7100
rect 20801 7098 20857 7100
rect 20561 7046 20607 7098
rect 20607 7046 20617 7098
rect 20641 7046 20671 7098
rect 20671 7046 20683 7098
rect 20683 7046 20697 7098
rect 20721 7046 20735 7098
rect 20735 7046 20747 7098
rect 20747 7046 20777 7098
rect 20801 7046 20811 7098
rect 20811 7046 20857 7098
rect 20561 7044 20617 7046
rect 20641 7044 20697 7046
rect 20721 7044 20777 7046
rect 20801 7044 20857 7046
rect 20561 6010 20617 6012
rect 20641 6010 20697 6012
rect 20721 6010 20777 6012
rect 20801 6010 20857 6012
rect 20561 5958 20607 6010
rect 20607 5958 20617 6010
rect 20641 5958 20671 6010
rect 20671 5958 20683 6010
rect 20683 5958 20697 6010
rect 20721 5958 20735 6010
rect 20735 5958 20747 6010
rect 20747 5958 20777 6010
rect 20801 5958 20811 6010
rect 20811 5958 20857 6010
rect 20561 5956 20617 5958
rect 20641 5956 20697 5958
rect 20721 5956 20777 5958
rect 20801 5956 20857 5958
rect 25134 17720 25190 17776
rect 24482 17434 24538 17436
rect 24562 17434 24618 17436
rect 24642 17434 24698 17436
rect 24722 17434 24778 17436
rect 24482 17382 24528 17434
rect 24528 17382 24538 17434
rect 24562 17382 24592 17434
rect 24592 17382 24604 17434
rect 24604 17382 24618 17434
rect 24642 17382 24656 17434
rect 24656 17382 24668 17434
rect 24668 17382 24698 17434
rect 24722 17382 24732 17434
rect 24732 17382 24778 17434
rect 24482 17380 24538 17382
rect 24562 17380 24618 17382
rect 24642 17380 24698 17382
rect 24722 17380 24778 17382
rect 25962 17856 26018 17912
rect 24214 15156 24270 15192
rect 24214 15136 24216 15156
rect 24216 15136 24268 15156
rect 24268 15136 24270 15156
rect 24482 16346 24538 16348
rect 24562 16346 24618 16348
rect 24642 16346 24698 16348
rect 24722 16346 24778 16348
rect 24482 16294 24528 16346
rect 24528 16294 24538 16346
rect 24562 16294 24592 16346
rect 24592 16294 24604 16346
rect 24604 16294 24618 16346
rect 24642 16294 24656 16346
rect 24656 16294 24668 16346
rect 24668 16294 24698 16346
rect 24722 16294 24732 16346
rect 24732 16294 24778 16346
rect 24482 16292 24538 16294
rect 24562 16292 24618 16294
rect 24642 16292 24698 16294
rect 24722 16292 24778 16294
rect 24482 15258 24538 15260
rect 24562 15258 24618 15260
rect 24642 15258 24698 15260
rect 24722 15258 24778 15260
rect 24482 15206 24528 15258
rect 24528 15206 24538 15258
rect 24562 15206 24592 15258
rect 24592 15206 24604 15258
rect 24604 15206 24618 15258
rect 24642 15206 24656 15258
rect 24656 15206 24668 15258
rect 24668 15206 24698 15258
rect 24722 15206 24732 15258
rect 24732 15206 24778 15258
rect 24482 15204 24538 15206
rect 24562 15204 24618 15206
rect 24642 15204 24698 15206
rect 24722 15204 24778 15206
rect 25870 15988 25872 16008
rect 25872 15988 25924 16008
rect 25924 15988 25926 16008
rect 25870 15952 25926 15988
rect 25410 15444 25412 15464
rect 25412 15444 25464 15464
rect 25464 15444 25466 15464
rect 25410 15408 25466 15444
rect 24482 14170 24538 14172
rect 24562 14170 24618 14172
rect 24642 14170 24698 14172
rect 24722 14170 24778 14172
rect 24482 14118 24528 14170
rect 24528 14118 24538 14170
rect 24562 14118 24592 14170
rect 24592 14118 24604 14170
rect 24604 14118 24618 14170
rect 24642 14118 24656 14170
rect 24656 14118 24668 14170
rect 24668 14118 24698 14170
rect 24722 14118 24732 14170
rect 24732 14118 24778 14170
rect 24482 14116 24538 14118
rect 24562 14116 24618 14118
rect 24642 14116 24698 14118
rect 24722 14116 24778 14118
rect 24214 13776 24270 13832
rect 24674 13252 24730 13288
rect 24674 13232 24676 13252
rect 24676 13232 24728 13252
rect 24728 13232 24730 13252
rect 24482 13082 24538 13084
rect 24562 13082 24618 13084
rect 24642 13082 24698 13084
rect 24722 13082 24778 13084
rect 24482 13030 24528 13082
rect 24528 13030 24538 13082
rect 24562 13030 24592 13082
rect 24592 13030 24604 13082
rect 24604 13030 24618 13082
rect 24642 13030 24656 13082
rect 24656 13030 24668 13082
rect 24668 13030 24698 13082
rect 24722 13030 24732 13082
rect 24732 13030 24778 13082
rect 24482 13028 24538 13030
rect 24562 13028 24618 13030
rect 24642 13028 24698 13030
rect 24722 13028 24778 13030
rect 24482 11994 24538 11996
rect 24562 11994 24618 11996
rect 24642 11994 24698 11996
rect 24722 11994 24778 11996
rect 24482 11942 24528 11994
rect 24528 11942 24538 11994
rect 24562 11942 24592 11994
rect 24592 11942 24604 11994
rect 24604 11942 24618 11994
rect 24642 11942 24656 11994
rect 24656 11942 24668 11994
rect 24668 11942 24698 11994
rect 24722 11942 24732 11994
rect 24732 11942 24778 11994
rect 24482 11940 24538 11942
rect 24562 11940 24618 11942
rect 24642 11940 24698 11942
rect 24722 11940 24778 11942
rect 28403 20154 28459 20156
rect 28483 20154 28539 20156
rect 28563 20154 28619 20156
rect 28643 20154 28699 20156
rect 28403 20102 28449 20154
rect 28449 20102 28459 20154
rect 28483 20102 28513 20154
rect 28513 20102 28525 20154
rect 28525 20102 28539 20154
rect 28563 20102 28577 20154
rect 28577 20102 28589 20154
rect 28589 20102 28619 20154
rect 28643 20102 28653 20154
rect 28653 20102 28699 20154
rect 28403 20100 28459 20102
rect 28483 20100 28539 20102
rect 28563 20100 28619 20102
rect 28643 20100 28699 20102
rect 28403 19066 28459 19068
rect 28483 19066 28539 19068
rect 28563 19066 28619 19068
rect 28643 19066 28699 19068
rect 28403 19014 28449 19066
rect 28449 19014 28459 19066
rect 28483 19014 28513 19066
rect 28513 19014 28525 19066
rect 28525 19014 28539 19066
rect 28563 19014 28577 19066
rect 28577 19014 28589 19066
rect 28589 19014 28619 19066
rect 28643 19014 28653 19066
rect 28653 19014 28699 19066
rect 28403 19012 28459 19014
rect 28483 19012 28539 19014
rect 28563 19012 28619 19014
rect 28643 19012 28699 19014
rect 26330 17584 26386 17640
rect 25962 14340 26018 14376
rect 25962 14320 25964 14340
rect 25964 14320 26016 14340
rect 26016 14320 26018 14340
rect 28403 17978 28459 17980
rect 28483 17978 28539 17980
rect 28563 17978 28619 17980
rect 28643 17978 28699 17980
rect 28403 17926 28449 17978
rect 28449 17926 28459 17978
rect 28483 17926 28513 17978
rect 28513 17926 28525 17978
rect 28525 17926 28539 17978
rect 28563 17926 28577 17978
rect 28577 17926 28589 17978
rect 28589 17926 28619 17978
rect 28643 17926 28653 17978
rect 28653 17926 28699 17978
rect 28403 17924 28459 17926
rect 28483 17924 28539 17926
rect 28563 17924 28619 17926
rect 28643 17924 28699 17926
rect 28403 16890 28459 16892
rect 28483 16890 28539 16892
rect 28563 16890 28619 16892
rect 28643 16890 28699 16892
rect 28403 16838 28449 16890
rect 28449 16838 28459 16890
rect 28483 16838 28513 16890
rect 28513 16838 28525 16890
rect 28525 16838 28539 16890
rect 28563 16838 28577 16890
rect 28577 16838 28589 16890
rect 28589 16838 28619 16890
rect 28643 16838 28653 16890
rect 28653 16838 28699 16890
rect 28403 16836 28459 16838
rect 28483 16836 28539 16838
rect 28563 16836 28619 16838
rect 28643 16836 28699 16838
rect 26422 15952 26478 16008
rect 26238 14456 26294 14512
rect 24482 10906 24538 10908
rect 24562 10906 24618 10908
rect 24642 10906 24698 10908
rect 24722 10906 24778 10908
rect 24482 10854 24528 10906
rect 24528 10854 24538 10906
rect 24562 10854 24592 10906
rect 24592 10854 24604 10906
rect 24604 10854 24618 10906
rect 24642 10854 24656 10906
rect 24656 10854 24668 10906
rect 24668 10854 24698 10906
rect 24722 10854 24732 10906
rect 24732 10854 24778 10906
rect 24482 10852 24538 10854
rect 24562 10852 24618 10854
rect 24642 10852 24698 10854
rect 24722 10852 24778 10854
rect 24482 9818 24538 9820
rect 24562 9818 24618 9820
rect 24642 9818 24698 9820
rect 24722 9818 24778 9820
rect 24482 9766 24528 9818
rect 24528 9766 24538 9818
rect 24562 9766 24592 9818
rect 24592 9766 24604 9818
rect 24604 9766 24618 9818
rect 24642 9766 24656 9818
rect 24656 9766 24668 9818
rect 24668 9766 24698 9818
rect 24722 9766 24732 9818
rect 24732 9766 24778 9818
rect 24482 9764 24538 9766
rect 24562 9764 24618 9766
rect 24642 9764 24698 9766
rect 24722 9764 24778 9766
rect 24482 8730 24538 8732
rect 24562 8730 24618 8732
rect 24642 8730 24698 8732
rect 24722 8730 24778 8732
rect 24482 8678 24528 8730
rect 24528 8678 24538 8730
rect 24562 8678 24592 8730
rect 24592 8678 24604 8730
rect 24604 8678 24618 8730
rect 24642 8678 24656 8730
rect 24656 8678 24668 8730
rect 24668 8678 24698 8730
rect 24722 8678 24732 8730
rect 24732 8678 24778 8730
rect 24482 8676 24538 8678
rect 24562 8676 24618 8678
rect 24642 8676 24698 8678
rect 24722 8676 24778 8678
rect 28403 15802 28459 15804
rect 28483 15802 28539 15804
rect 28563 15802 28619 15804
rect 28643 15802 28699 15804
rect 28403 15750 28449 15802
rect 28449 15750 28459 15802
rect 28483 15750 28513 15802
rect 28513 15750 28525 15802
rect 28525 15750 28539 15802
rect 28563 15750 28577 15802
rect 28577 15750 28589 15802
rect 28589 15750 28619 15802
rect 28643 15750 28653 15802
rect 28653 15750 28699 15802
rect 28403 15748 28459 15750
rect 28483 15748 28539 15750
rect 28563 15748 28619 15750
rect 28643 15748 28699 15750
rect 25410 9016 25466 9072
rect 28403 14714 28459 14716
rect 28483 14714 28539 14716
rect 28563 14714 28619 14716
rect 28643 14714 28699 14716
rect 28403 14662 28449 14714
rect 28449 14662 28459 14714
rect 28483 14662 28513 14714
rect 28513 14662 28525 14714
rect 28525 14662 28539 14714
rect 28563 14662 28577 14714
rect 28577 14662 28589 14714
rect 28589 14662 28619 14714
rect 28643 14662 28653 14714
rect 28653 14662 28699 14714
rect 28403 14660 28459 14662
rect 28483 14660 28539 14662
rect 28563 14660 28619 14662
rect 28643 14660 28699 14662
rect 28722 14456 28778 14512
rect 28814 14340 28870 14376
rect 28814 14320 28816 14340
rect 28816 14320 28868 14340
rect 28868 14320 28870 14340
rect 28403 13626 28459 13628
rect 28483 13626 28539 13628
rect 28563 13626 28619 13628
rect 28643 13626 28699 13628
rect 28403 13574 28449 13626
rect 28449 13574 28459 13626
rect 28483 13574 28513 13626
rect 28513 13574 28525 13626
rect 28525 13574 28539 13626
rect 28563 13574 28577 13626
rect 28577 13574 28589 13626
rect 28589 13574 28619 13626
rect 28643 13574 28653 13626
rect 28653 13574 28699 13626
rect 28403 13572 28459 13574
rect 28483 13572 28539 13574
rect 28563 13572 28619 13574
rect 28643 13572 28699 13574
rect 28403 12538 28459 12540
rect 28483 12538 28539 12540
rect 28563 12538 28619 12540
rect 28643 12538 28699 12540
rect 28403 12486 28449 12538
rect 28449 12486 28459 12538
rect 28483 12486 28513 12538
rect 28513 12486 28525 12538
rect 28525 12486 28539 12538
rect 28563 12486 28577 12538
rect 28577 12486 28589 12538
rect 28589 12486 28619 12538
rect 28643 12486 28653 12538
rect 28653 12486 28699 12538
rect 28403 12484 28459 12486
rect 28483 12484 28539 12486
rect 28563 12484 28619 12486
rect 28643 12484 28699 12486
rect 28403 11450 28459 11452
rect 28483 11450 28539 11452
rect 28563 11450 28619 11452
rect 28643 11450 28699 11452
rect 28403 11398 28449 11450
rect 28449 11398 28459 11450
rect 28483 11398 28513 11450
rect 28513 11398 28525 11450
rect 28525 11398 28539 11450
rect 28563 11398 28577 11450
rect 28577 11398 28589 11450
rect 28589 11398 28619 11450
rect 28643 11398 28653 11450
rect 28653 11398 28699 11450
rect 28403 11396 28459 11398
rect 28483 11396 28539 11398
rect 28563 11396 28619 11398
rect 28643 11396 28699 11398
rect 26974 9016 27030 9072
rect 28403 10362 28459 10364
rect 28483 10362 28539 10364
rect 28563 10362 28619 10364
rect 28643 10362 28699 10364
rect 28403 10310 28449 10362
rect 28449 10310 28459 10362
rect 28483 10310 28513 10362
rect 28513 10310 28525 10362
rect 28525 10310 28539 10362
rect 28563 10310 28577 10362
rect 28577 10310 28589 10362
rect 28589 10310 28619 10362
rect 28643 10310 28653 10362
rect 28653 10310 28699 10362
rect 28403 10308 28459 10310
rect 28483 10308 28539 10310
rect 28563 10308 28619 10310
rect 28643 10308 28699 10310
rect 28403 9274 28459 9276
rect 28483 9274 28539 9276
rect 28563 9274 28619 9276
rect 28643 9274 28699 9276
rect 28403 9222 28449 9274
rect 28449 9222 28459 9274
rect 28483 9222 28513 9274
rect 28513 9222 28525 9274
rect 28525 9222 28539 9274
rect 28563 9222 28577 9274
rect 28577 9222 28589 9274
rect 28589 9222 28619 9274
rect 28643 9222 28653 9274
rect 28653 9222 28699 9274
rect 28403 9220 28459 9222
rect 28483 9220 28539 9222
rect 28563 9220 28619 9222
rect 28643 9220 28699 9222
rect 30286 16904 30342 16960
rect 31758 17856 31814 17912
rect 32324 20698 32380 20700
rect 32404 20698 32460 20700
rect 32484 20698 32540 20700
rect 32564 20698 32620 20700
rect 32324 20646 32370 20698
rect 32370 20646 32380 20698
rect 32404 20646 32434 20698
rect 32434 20646 32446 20698
rect 32446 20646 32460 20698
rect 32484 20646 32498 20698
rect 32498 20646 32510 20698
rect 32510 20646 32540 20698
rect 32564 20646 32574 20698
rect 32574 20646 32620 20698
rect 32324 20644 32380 20646
rect 32404 20644 32460 20646
rect 32484 20644 32540 20646
rect 32564 20644 32620 20646
rect 32324 19610 32380 19612
rect 32404 19610 32460 19612
rect 32484 19610 32540 19612
rect 32564 19610 32620 19612
rect 32324 19558 32370 19610
rect 32370 19558 32380 19610
rect 32404 19558 32434 19610
rect 32434 19558 32446 19610
rect 32446 19558 32460 19610
rect 32484 19558 32498 19610
rect 32498 19558 32510 19610
rect 32510 19558 32540 19610
rect 32564 19558 32574 19610
rect 32574 19558 32620 19610
rect 32324 19556 32380 19558
rect 32404 19556 32460 19558
rect 32484 19556 32540 19558
rect 32564 19556 32620 19558
rect 32324 18522 32380 18524
rect 32404 18522 32460 18524
rect 32484 18522 32540 18524
rect 32564 18522 32620 18524
rect 32324 18470 32370 18522
rect 32370 18470 32380 18522
rect 32404 18470 32434 18522
rect 32434 18470 32446 18522
rect 32446 18470 32460 18522
rect 32484 18470 32498 18522
rect 32498 18470 32510 18522
rect 32510 18470 32540 18522
rect 32564 18470 32574 18522
rect 32574 18470 32620 18522
rect 32324 18468 32380 18470
rect 32404 18468 32460 18470
rect 32484 18468 32540 18470
rect 32564 18468 32620 18470
rect 32324 17434 32380 17436
rect 32404 17434 32460 17436
rect 32484 17434 32540 17436
rect 32564 17434 32620 17436
rect 32324 17382 32370 17434
rect 32370 17382 32380 17434
rect 32404 17382 32434 17434
rect 32434 17382 32446 17434
rect 32446 17382 32460 17434
rect 32484 17382 32498 17434
rect 32498 17382 32510 17434
rect 32510 17382 32540 17434
rect 32564 17382 32574 17434
rect 32574 17382 32620 17434
rect 32324 17380 32380 17382
rect 32404 17380 32460 17382
rect 32484 17380 32540 17382
rect 32564 17380 32620 17382
rect 32324 16346 32380 16348
rect 32404 16346 32460 16348
rect 32484 16346 32540 16348
rect 32564 16346 32620 16348
rect 32324 16294 32370 16346
rect 32370 16294 32380 16346
rect 32404 16294 32434 16346
rect 32434 16294 32446 16346
rect 32446 16294 32460 16346
rect 32484 16294 32498 16346
rect 32498 16294 32510 16346
rect 32510 16294 32540 16346
rect 32564 16294 32574 16346
rect 32574 16294 32620 16346
rect 32324 16292 32380 16294
rect 32404 16292 32460 16294
rect 32484 16292 32540 16294
rect 32564 16292 32620 16294
rect 32324 15258 32380 15260
rect 32404 15258 32460 15260
rect 32484 15258 32540 15260
rect 32564 15258 32620 15260
rect 32324 15206 32370 15258
rect 32370 15206 32380 15258
rect 32404 15206 32434 15258
rect 32434 15206 32446 15258
rect 32446 15206 32460 15258
rect 32484 15206 32498 15258
rect 32498 15206 32510 15258
rect 32510 15206 32540 15258
rect 32564 15206 32574 15258
rect 32574 15206 32620 15258
rect 32324 15204 32380 15206
rect 32404 15204 32460 15206
rect 32484 15204 32540 15206
rect 32564 15204 32620 15206
rect 32324 14170 32380 14172
rect 32404 14170 32460 14172
rect 32484 14170 32540 14172
rect 32564 14170 32620 14172
rect 32324 14118 32370 14170
rect 32370 14118 32380 14170
rect 32404 14118 32434 14170
rect 32434 14118 32446 14170
rect 32446 14118 32460 14170
rect 32484 14118 32498 14170
rect 32498 14118 32510 14170
rect 32510 14118 32540 14170
rect 32564 14118 32574 14170
rect 32574 14118 32620 14170
rect 32324 14116 32380 14118
rect 32404 14116 32460 14118
rect 32484 14116 32540 14118
rect 32564 14116 32620 14118
rect 32324 13082 32380 13084
rect 32404 13082 32460 13084
rect 32484 13082 32540 13084
rect 32564 13082 32620 13084
rect 32324 13030 32370 13082
rect 32370 13030 32380 13082
rect 32404 13030 32434 13082
rect 32434 13030 32446 13082
rect 32446 13030 32460 13082
rect 32484 13030 32498 13082
rect 32498 13030 32510 13082
rect 32510 13030 32540 13082
rect 32564 13030 32574 13082
rect 32574 13030 32620 13082
rect 32324 13028 32380 13030
rect 32404 13028 32460 13030
rect 32484 13028 32540 13030
rect 32564 13028 32620 13030
rect 32324 11994 32380 11996
rect 32404 11994 32460 11996
rect 32484 11994 32540 11996
rect 32564 11994 32620 11996
rect 32324 11942 32370 11994
rect 32370 11942 32380 11994
rect 32404 11942 32434 11994
rect 32434 11942 32446 11994
rect 32446 11942 32460 11994
rect 32484 11942 32498 11994
rect 32498 11942 32510 11994
rect 32510 11942 32540 11994
rect 32564 11942 32574 11994
rect 32574 11942 32620 11994
rect 32324 11940 32380 11942
rect 32404 11940 32460 11942
rect 32484 11940 32540 11942
rect 32564 11940 32620 11942
rect 32324 10906 32380 10908
rect 32404 10906 32460 10908
rect 32484 10906 32540 10908
rect 32564 10906 32620 10908
rect 32324 10854 32370 10906
rect 32370 10854 32380 10906
rect 32404 10854 32434 10906
rect 32434 10854 32446 10906
rect 32446 10854 32460 10906
rect 32484 10854 32498 10906
rect 32498 10854 32510 10906
rect 32510 10854 32540 10906
rect 32564 10854 32574 10906
rect 32574 10854 32620 10906
rect 32324 10852 32380 10854
rect 32404 10852 32460 10854
rect 32484 10852 32540 10854
rect 32564 10852 32620 10854
rect 32324 9818 32380 9820
rect 32404 9818 32460 9820
rect 32484 9818 32540 9820
rect 32564 9818 32620 9820
rect 32324 9766 32370 9818
rect 32370 9766 32380 9818
rect 32404 9766 32434 9818
rect 32434 9766 32446 9818
rect 32446 9766 32460 9818
rect 32484 9766 32498 9818
rect 32498 9766 32510 9818
rect 32510 9766 32540 9818
rect 32564 9766 32574 9818
rect 32574 9766 32620 9818
rect 32324 9764 32380 9766
rect 32404 9764 32460 9766
rect 32484 9764 32540 9766
rect 32564 9764 32620 9766
rect 32324 8730 32380 8732
rect 32404 8730 32460 8732
rect 32484 8730 32540 8732
rect 32564 8730 32620 8732
rect 32324 8678 32370 8730
rect 32370 8678 32380 8730
rect 32404 8678 32434 8730
rect 32434 8678 32446 8730
rect 32446 8678 32460 8730
rect 32484 8678 32498 8730
rect 32498 8678 32510 8730
rect 32510 8678 32540 8730
rect 32564 8678 32574 8730
rect 32574 8678 32620 8730
rect 32324 8676 32380 8678
rect 32404 8676 32460 8678
rect 32484 8676 32540 8678
rect 32564 8676 32620 8678
rect 28403 8186 28459 8188
rect 28483 8186 28539 8188
rect 28563 8186 28619 8188
rect 28643 8186 28699 8188
rect 28403 8134 28449 8186
rect 28449 8134 28459 8186
rect 28483 8134 28513 8186
rect 28513 8134 28525 8186
rect 28525 8134 28539 8186
rect 28563 8134 28577 8186
rect 28577 8134 28589 8186
rect 28589 8134 28619 8186
rect 28643 8134 28653 8186
rect 28653 8134 28699 8186
rect 28403 8132 28459 8134
rect 28483 8132 28539 8134
rect 28563 8132 28619 8134
rect 28643 8132 28699 8134
rect 24482 7642 24538 7644
rect 24562 7642 24618 7644
rect 24642 7642 24698 7644
rect 24722 7642 24778 7644
rect 24482 7590 24528 7642
rect 24528 7590 24538 7642
rect 24562 7590 24592 7642
rect 24592 7590 24604 7642
rect 24604 7590 24618 7642
rect 24642 7590 24656 7642
rect 24656 7590 24668 7642
rect 24668 7590 24698 7642
rect 24722 7590 24732 7642
rect 24732 7590 24778 7642
rect 24482 7588 24538 7590
rect 24562 7588 24618 7590
rect 24642 7588 24698 7590
rect 24722 7588 24778 7590
rect 32324 7642 32380 7644
rect 32404 7642 32460 7644
rect 32484 7642 32540 7644
rect 32564 7642 32620 7644
rect 32324 7590 32370 7642
rect 32370 7590 32380 7642
rect 32404 7590 32434 7642
rect 32434 7590 32446 7642
rect 32446 7590 32460 7642
rect 32484 7590 32498 7642
rect 32498 7590 32510 7642
rect 32510 7590 32540 7642
rect 32564 7590 32574 7642
rect 32574 7590 32620 7642
rect 32324 7588 32380 7590
rect 32404 7588 32460 7590
rect 32484 7588 32540 7590
rect 32564 7588 32620 7590
rect 28403 7098 28459 7100
rect 28483 7098 28539 7100
rect 28563 7098 28619 7100
rect 28643 7098 28699 7100
rect 28403 7046 28449 7098
rect 28449 7046 28459 7098
rect 28483 7046 28513 7098
rect 28513 7046 28525 7098
rect 28525 7046 28539 7098
rect 28563 7046 28577 7098
rect 28577 7046 28589 7098
rect 28589 7046 28619 7098
rect 28643 7046 28653 7098
rect 28653 7046 28699 7098
rect 28403 7044 28459 7046
rect 28483 7044 28539 7046
rect 28563 7044 28619 7046
rect 28643 7044 28699 7046
rect 24482 6554 24538 6556
rect 24562 6554 24618 6556
rect 24642 6554 24698 6556
rect 24722 6554 24778 6556
rect 24482 6502 24528 6554
rect 24528 6502 24538 6554
rect 24562 6502 24592 6554
rect 24592 6502 24604 6554
rect 24604 6502 24618 6554
rect 24642 6502 24656 6554
rect 24656 6502 24668 6554
rect 24668 6502 24698 6554
rect 24722 6502 24732 6554
rect 24732 6502 24778 6554
rect 24482 6500 24538 6502
rect 24562 6500 24618 6502
rect 24642 6500 24698 6502
rect 24722 6500 24778 6502
rect 32324 6554 32380 6556
rect 32404 6554 32460 6556
rect 32484 6554 32540 6556
rect 32564 6554 32620 6556
rect 32324 6502 32370 6554
rect 32370 6502 32380 6554
rect 32404 6502 32434 6554
rect 32434 6502 32446 6554
rect 32446 6502 32460 6554
rect 32484 6502 32498 6554
rect 32498 6502 32510 6554
rect 32510 6502 32540 6554
rect 32564 6502 32574 6554
rect 32574 6502 32620 6554
rect 32324 6500 32380 6502
rect 32404 6500 32460 6502
rect 32484 6500 32540 6502
rect 32564 6500 32620 6502
rect 28403 6010 28459 6012
rect 28483 6010 28539 6012
rect 28563 6010 28619 6012
rect 28643 6010 28699 6012
rect 28403 5958 28449 6010
rect 28449 5958 28459 6010
rect 28483 5958 28513 6010
rect 28513 5958 28525 6010
rect 28525 5958 28539 6010
rect 28563 5958 28577 6010
rect 28577 5958 28589 6010
rect 28589 5958 28619 6010
rect 28643 5958 28653 6010
rect 28653 5958 28699 6010
rect 28403 5956 28459 5958
rect 28483 5956 28539 5958
rect 28563 5956 28619 5958
rect 28643 5956 28699 5958
rect 24482 5466 24538 5468
rect 24562 5466 24618 5468
rect 24642 5466 24698 5468
rect 24722 5466 24778 5468
rect 24482 5414 24528 5466
rect 24528 5414 24538 5466
rect 24562 5414 24592 5466
rect 24592 5414 24604 5466
rect 24604 5414 24618 5466
rect 24642 5414 24656 5466
rect 24656 5414 24668 5466
rect 24668 5414 24698 5466
rect 24722 5414 24732 5466
rect 24732 5414 24778 5466
rect 24482 5412 24538 5414
rect 24562 5412 24618 5414
rect 24642 5412 24698 5414
rect 24722 5412 24778 5414
rect 32324 5466 32380 5468
rect 32404 5466 32460 5468
rect 32484 5466 32540 5468
rect 32564 5466 32620 5468
rect 32324 5414 32370 5466
rect 32370 5414 32380 5466
rect 32404 5414 32434 5466
rect 32434 5414 32446 5466
rect 32446 5414 32460 5466
rect 32484 5414 32498 5466
rect 32498 5414 32510 5466
rect 32510 5414 32540 5466
rect 32564 5414 32574 5466
rect 32574 5414 32620 5466
rect 32324 5412 32380 5414
rect 32404 5412 32460 5414
rect 32484 5412 32540 5414
rect 32564 5412 32620 5414
rect 4877 4922 4933 4924
rect 4957 4922 5013 4924
rect 5037 4922 5093 4924
rect 5117 4922 5173 4924
rect 4877 4870 4923 4922
rect 4923 4870 4933 4922
rect 4957 4870 4987 4922
rect 4987 4870 4999 4922
rect 4999 4870 5013 4922
rect 5037 4870 5051 4922
rect 5051 4870 5063 4922
rect 5063 4870 5093 4922
rect 5117 4870 5127 4922
rect 5127 4870 5173 4922
rect 4877 4868 4933 4870
rect 4957 4868 5013 4870
rect 5037 4868 5093 4870
rect 5117 4868 5173 4870
rect 12719 4922 12775 4924
rect 12799 4922 12855 4924
rect 12879 4922 12935 4924
rect 12959 4922 13015 4924
rect 12719 4870 12765 4922
rect 12765 4870 12775 4922
rect 12799 4870 12829 4922
rect 12829 4870 12841 4922
rect 12841 4870 12855 4922
rect 12879 4870 12893 4922
rect 12893 4870 12905 4922
rect 12905 4870 12935 4922
rect 12959 4870 12969 4922
rect 12969 4870 13015 4922
rect 12719 4868 12775 4870
rect 12799 4868 12855 4870
rect 12879 4868 12935 4870
rect 12959 4868 13015 4870
rect 20561 4922 20617 4924
rect 20641 4922 20697 4924
rect 20721 4922 20777 4924
rect 20801 4922 20857 4924
rect 20561 4870 20607 4922
rect 20607 4870 20617 4922
rect 20641 4870 20671 4922
rect 20671 4870 20683 4922
rect 20683 4870 20697 4922
rect 20721 4870 20735 4922
rect 20735 4870 20747 4922
rect 20747 4870 20777 4922
rect 20801 4870 20811 4922
rect 20811 4870 20857 4922
rect 20561 4868 20617 4870
rect 20641 4868 20697 4870
rect 20721 4868 20777 4870
rect 20801 4868 20857 4870
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28643 4922 28699 4924
rect 28403 4870 28449 4922
rect 28449 4870 28459 4922
rect 28483 4870 28513 4922
rect 28513 4870 28525 4922
rect 28525 4870 28539 4922
rect 28563 4870 28577 4922
rect 28577 4870 28589 4922
rect 28589 4870 28619 4922
rect 28643 4870 28653 4922
rect 28653 4870 28699 4922
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 28643 4868 28699 4870
rect 8798 4378 8854 4380
rect 8878 4378 8934 4380
rect 8958 4378 9014 4380
rect 9038 4378 9094 4380
rect 8798 4326 8844 4378
rect 8844 4326 8854 4378
rect 8878 4326 8908 4378
rect 8908 4326 8920 4378
rect 8920 4326 8934 4378
rect 8958 4326 8972 4378
rect 8972 4326 8984 4378
rect 8984 4326 9014 4378
rect 9038 4326 9048 4378
rect 9048 4326 9094 4378
rect 8798 4324 8854 4326
rect 8878 4324 8934 4326
rect 8958 4324 9014 4326
rect 9038 4324 9094 4326
rect 16640 4378 16696 4380
rect 16720 4378 16776 4380
rect 16800 4378 16856 4380
rect 16880 4378 16936 4380
rect 16640 4326 16686 4378
rect 16686 4326 16696 4378
rect 16720 4326 16750 4378
rect 16750 4326 16762 4378
rect 16762 4326 16776 4378
rect 16800 4326 16814 4378
rect 16814 4326 16826 4378
rect 16826 4326 16856 4378
rect 16880 4326 16890 4378
rect 16890 4326 16936 4378
rect 16640 4324 16696 4326
rect 16720 4324 16776 4326
rect 16800 4324 16856 4326
rect 16880 4324 16936 4326
rect 24482 4378 24538 4380
rect 24562 4378 24618 4380
rect 24642 4378 24698 4380
rect 24722 4378 24778 4380
rect 24482 4326 24528 4378
rect 24528 4326 24538 4378
rect 24562 4326 24592 4378
rect 24592 4326 24604 4378
rect 24604 4326 24618 4378
rect 24642 4326 24656 4378
rect 24656 4326 24668 4378
rect 24668 4326 24698 4378
rect 24722 4326 24732 4378
rect 24732 4326 24778 4378
rect 24482 4324 24538 4326
rect 24562 4324 24618 4326
rect 24642 4324 24698 4326
rect 24722 4324 24778 4326
rect 32324 4378 32380 4380
rect 32404 4378 32460 4380
rect 32484 4378 32540 4380
rect 32564 4378 32620 4380
rect 32324 4326 32370 4378
rect 32370 4326 32380 4378
rect 32404 4326 32434 4378
rect 32434 4326 32446 4378
rect 32446 4326 32460 4378
rect 32484 4326 32498 4378
rect 32498 4326 32510 4378
rect 32510 4326 32540 4378
rect 32564 4326 32574 4378
rect 32574 4326 32620 4378
rect 32324 4324 32380 4326
rect 32404 4324 32460 4326
rect 32484 4324 32540 4326
rect 32564 4324 32620 4326
rect 4877 3834 4933 3836
rect 4957 3834 5013 3836
rect 5037 3834 5093 3836
rect 5117 3834 5173 3836
rect 4877 3782 4923 3834
rect 4923 3782 4933 3834
rect 4957 3782 4987 3834
rect 4987 3782 4999 3834
rect 4999 3782 5013 3834
rect 5037 3782 5051 3834
rect 5051 3782 5063 3834
rect 5063 3782 5093 3834
rect 5117 3782 5127 3834
rect 5127 3782 5173 3834
rect 4877 3780 4933 3782
rect 4957 3780 5013 3782
rect 5037 3780 5093 3782
rect 5117 3780 5173 3782
rect 12719 3834 12775 3836
rect 12799 3834 12855 3836
rect 12879 3834 12935 3836
rect 12959 3834 13015 3836
rect 12719 3782 12765 3834
rect 12765 3782 12775 3834
rect 12799 3782 12829 3834
rect 12829 3782 12841 3834
rect 12841 3782 12855 3834
rect 12879 3782 12893 3834
rect 12893 3782 12905 3834
rect 12905 3782 12935 3834
rect 12959 3782 12969 3834
rect 12969 3782 13015 3834
rect 12719 3780 12775 3782
rect 12799 3780 12855 3782
rect 12879 3780 12935 3782
rect 12959 3780 13015 3782
rect 20561 3834 20617 3836
rect 20641 3834 20697 3836
rect 20721 3834 20777 3836
rect 20801 3834 20857 3836
rect 20561 3782 20607 3834
rect 20607 3782 20617 3834
rect 20641 3782 20671 3834
rect 20671 3782 20683 3834
rect 20683 3782 20697 3834
rect 20721 3782 20735 3834
rect 20735 3782 20747 3834
rect 20747 3782 20777 3834
rect 20801 3782 20811 3834
rect 20811 3782 20857 3834
rect 20561 3780 20617 3782
rect 20641 3780 20697 3782
rect 20721 3780 20777 3782
rect 20801 3780 20857 3782
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28643 3834 28699 3836
rect 28403 3782 28449 3834
rect 28449 3782 28459 3834
rect 28483 3782 28513 3834
rect 28513 3782 28525 3834
rect 28525 3782 28539 3834
rect 28563 3782 28577 3834
rect 28577 3782 28589 3834
rect 28589 3782 28619 3834
rect 28643 3782 28653 3834
rect 28653 3782 28699 3834
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28643 3780 28699 3782
rect 8798 3290 8854 3292
rect 8878 3290 8934 3292
rect 8958 3290 9014 3292
rect 9038 3290 9094 3292
rect 8798 3238 8844 3290
rect 8844 3238 8854 3290
rect 8878 3238 8908 3290
rect 8908 3238 8920 3290
rect 8920 3238 8934 3290
rect 8958 3238 8972 3290
rect 8972 3238 8984 3290
rect 8984 3238 9014 3290
rect 9038 3238 9048 3290
rect 9048 3238 9094 3290
rect 8798 3236 8854 3238
rect 8878 3236 8934 3238
rect 8958 3236 9014 3238
rect 9038 3236 9094 3238
rect 16640 3290 16696 3292
rect 16720 3290 16776 3292
rect 16800 3290 16856 3292
rect 16880 3290 16936 3292
rect 16640 3238 16686 3290
rect 16686 3238 16696 3290
rect 16720 3238 16750 3290
rect 16750 3238 16762 3290
rect 16762 3238 16776 3290
rect 16800 3238 16814 3290
rect 16814 3238 16826 3290
rect 16826 3238 16856 3290
rect 16880 3238 16890 3290
rect 16890 3238 16936 3290
rect 16640 3236 16696 3238
rect 16720 3236 16776 3238
rect 16800 3236 16856 3238
rect 16880 3236 16936 3238
rect 24482 3290 24538 3292
rect 24562 3290 24618 3292
rect 24642 3290 24698 3292
rect 24722 3290 24778 3292
rect 24482 3238 24528 3290
rect 24528 3238 24538 3290
rect 24562 3238 24592 3290
rect 24592 3238 24604 3290
rect 24604 3238 24618 3290
rect 24642 3238 24656 3290
rect 24656 3238 24668 3290
rect 24668 3238 24698 3290
rect 24722 3238 24732 3290
rect 24732 3238 24778 3290
rect 24482 3236 24538 3238
rect 24562 3236 24618 3238
rect 24642 3236 24698 3238
rect 24722 3236 24778 3238
rect 32324 3290 32380 3292
rect 32404 3290 32460 3292
rect 32484 3290 32540 3292
rect 32564 3290 32620 3292
rect 32324 3238 32370 3290
rect 32370 3238 32380 3290
rect 32404 3238 32434 3290
rect 32434 3238 32446 3290
rect 32446 3238 32460 3290
rect 32484 3238 32498 3290
rect 32498 3238 32510 3290
rect 32510 3238 32540 3290
rect 32564 3238 32574 3290
rect 32574 3238 32620 3290
rect 32324 3236 32380 3238
rect 32404 3236 32460 3238
rect 32484 3236 32540 3238
rect 32564 3236 32620 3238
rect 4877 2746 4933 2748
rect 4957 2746 5013 2748
rect 5037 2746 5093 2748
rect 5117 2746 5173 2748
rect 4877 2694 4923 2746
rect 4923 2694 4933 2746
rect 4957 2694 4987 2746
rect 4987 2694 4999 2746
rect 4999 2694 5013 2746
rect 5037 2694 5051 2746
rect 5051 2694 5063 2746
rect 5063 2694 5093 2746
rect 5117 2694 5127 2746
rect 5127 2694 5173 2746
rect 4877 2692 4933 2694
rect 4957 2692 5013 2694
rect 5037 2692 5093 2694
rect 5117 2692 5173 2694
rect 12719 2746 12775 2748
rect 12799 2746 12855 2748
rect 12879 2746 12935 2748
rect 12959 2746 13015 2748
rect 12719 2694 12765 2746
rect 12765 2694 12775 2746
rect 12799 2694 12829 2746
rect 12829 2694 12841 2746
rect 12841 2694 12855 2746
rect 12879 2694 12893 2746
rect 12893 2694 12905 2746
rect 12905 2694 12935 2746
rect 12959 2694 12969 2746
rect 12969 2694 13015 2746
rect 12719 2692 12775 2694
rect 12799 2692 12855 2694
rect 12879 2692 12935 2694
rect 12959 2692 13015 2694
rect 20561 2746 20617 2748
rect 20641 2746 20697 2748
rect 20721 2746 20777 2748
rect 20801 2746 20857 2748
rect 20561 2694 20607 2746
rect 20607 2694 20617 2746
rect 20641 2694 20671 2746
rect 20671 2694 20683 2746
rect 20683 2694 20697 2746
rect 20721 2694 20735 2746
rect 20735 2694 20747 2746
rect 20747 2694 20777 2746
rect 20801 2694 20811 2746
rect 20811 2694 20857 2746
rect 20561 2692 20617 2694
rect 20641 2692 20697 2694
rect 20721 2692 20777 2694
rect 20801 2692 20857 2694
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28643 2746 28699 2748
rect 28403 2694 28449 2746
rect 28449 2694 28459 2746
rect 28483 2694 28513 2746
rect 28513 2694 28525 2746
rect 28525 2694 28539 2746
rect 28563 2694 28577 2746
rect 28577 2694 28589 2746
rect 28589 2694 28619 2746
rect 28643 2694 28653 2746
rect 28653 2694 28699 2746
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 28643 2692 28699 2694
rect 8798 2202 8854 2204
rect 8878 2202 8934 2204
rect 8958 2202 9014 2204
rect 9038 2202 9094 2204
rect 8798 2150 8844 2202
rect 8844 2150 8854 2202
rect 8878 2150 8908 2202
rect 8908 2150 8920 2202
rect 8920 2150 8934 2202
rect 8958 2150 8972 2202
rect 8972 2150 8984 2202
rect 8984 2150 9014 2202
rect 9038 2150 9048 2202
rect 9048 2150 9094 2202
rect 8798 2148 8854 2150
rect 8878 2148 8934 2150
rect 8958 2148 9014 2150
rect 9038 2148 9094 2150
rect 16640 2202 16696 2204
rect 16720 2202 16776 2204
rect 16800 2202 16856 2204
rect 16880 2202 16936 2204
rect 16640 2150 16686 2202
rect 16686 2150 16696 2202
rect 16720 2150 16750 2202
rect 16750 2150 16762 2202
rect 16762 2150 16776 2202
rect 16800 2150 16814 2202
rect 16814 2150 16826 2202
rect 16826 2150 16856 2202
rect 16880 2150 16890 2202
rect 16890 2150 16936 2202
rect 16640 2148 16696 2150
rect 16720 2148 16776 2150
rect 16800 2148 16856 2150
rect 16880 2148 16936 2150
rect 24482 2202 24538 2204
rect 24562 2202 24618 2204
rect 24642 2202 24698 2204
rect 24722 2202 24778 2204
rect 24482 2150 24528 2202
rect 24528 2150 24538 2202
rect 24562 2150 24592 2202
rect 24592 2150 24604 2202
rect 24604 2150 24618 2202
rect 24642 2150 24656 2202
rect 24656 2150 24668 2202
rect 24668 2150 24698 2202
rect 24722 2150 24732 2202
rect 24732 2150 24778 2202
rect 24482 2148 24538 2150
rect 24562 2148 24618 2150
rect 24642 2148 24698 2150
rect 24722 2148 24778 2150
rect 32324 2202 32380 2204
rect 32404 2202 32460 2204
rect 32484 2202 32540 2204
rect 32564 2202 32620 2204
rect 32324 2150 32370 2202
rect 32370 2150 32380 2202
rect 32404 2150 32434 2202
rect 32434 2150 32446 2202
rect 32446 2150 32460 2202
rect 32484 2150 32498 2202
rect 32498 2150 32510 2202
rect 32510 2150 32540 2202
rect 32564 2150 32574 2202
rect 32574 2150 32620 2202
rect 32324 2148 32380 2150
rect 32404 2148 32460 2150
rect 32484 2148 32540 2150
rect 32564 2148 32620 2150
rect 4877 1658 4933 1660
rect 4957 1658 5013 1660
rect 5037 1658 5093 1660
rect 5117 1658 5173 1660
rect 4877 1606 4923 1658
rect 4923 1606 4933 1658
rect 4957 1606 4987 1658
rect 4987 1606 4999 1658
rect 4999 1606 5013 1658
rect 5037 1606 5051 1658
rect 5051 1606 5063 1658
rect 5063 1606 5093 1658
rect 5117 1606 5127 1658
rect 5127 1606 5173 1658
rect 4877 1604 4933 1606
rect 4957 1604 5013 1606
rect 5037 1604 5093 1606
rect 5117 1604 5173 1606
rect 12719 1658 12775 1660
rect 12799 1658 12855 1660
rect 12879 1658 12935 1660
rect 12959 1658 13015 1660
rect 12719 1606 12765 1658
rect 12765 1606 12775 1658
rect 12799 1606 12829 1658
rect 12829 1606 12841 1658
rect 12841 1606 12855 1658
rect 12879 1606 12893 1658
rect 12893 1606 12905 1658
rect 12905 1606 12935 1658
rect 12959 1606 12969 1658
rect 12969 1606 13015 1658
rect 12719 1604 12775 1606
rect 12799 1604 12855 1606
rect 12879 1604 12935 1606
rect 12959 1604 13015 1606
rect 20561 1658 20617 1660
rect 20641 1658 20697 1660
rect 20721 1658 20777 1660
rect 20801 1658 20857 1660
rect 20561 1606 20607 1658
rect 20607 1606 20617 1658
rect 20641 1606 20671 1658
rect 20671 1606 20683 1658
rect 20683 1606 20697 1658
rect 20721 1606 20735 1658
rect 20735 1606 20747 1658
rect 20747 1606 20777 1658
rect 20801 1606 20811 1658
rect 20811 1606 20857 1658
rect 20561 1604 20617 1606
rect 20641 1604 20697 1606
rect 20721 1604 20777 1606
rect 20801 1604 20857 1606
rect 28403 1658 28459 1660
rect 28483 1658 28539 1660
rect 28563 1658 28619 1660
rect 28643 1658 28699 1660
rect 28403 1606 28449 1658
rect 28449 1606 28459 1658
rect 28483 1606 28513 1658
rect 28513 1606 28525 1658
rect 28525 1606 28539 1658
rect 28563 1606 28577 1658
rect 28577 1606 28589 1658
rect 28589 1606 28619 1658
rect 28643 1606 28653 1658
rect 28653 1606 28699 1658
rect 28403 1604 28459 1606
rect 28483 1604 28539 1606
rect 28563 1604 28619 1606
rect 28643 1604 28699 1606
rect 8798 1114 8854 1116
rect 8878 1114 8934 1116
rect 8958 1114 9014 1116
rect 9038 1114 9094 1116
rect 8798 1062 8844 1114
rect 8844 1062 8854 1114
rect 8878 1062 8908 1114
rect 8908 1062 8920 1114
rect 8920 1062 8934 1114
rect 8958 1062 8972 1114
rect 8972 1062 8984 1114
rect 8984 1062 9014 1114
rect 9038 1062 9048 1114
rect 9048 1062 9094 1114
rect 8798 1060 8854 1062
rect 8878 1060 8934 1062
rect 8958 1060 9014 1062
rect 9038 1060 9094 1062
rect 16640 1114 16696 1116
rect 16720 1114 16776 1116
rect 16800 1114 16856 1116
rect 16880 1114 16936 1116
rect 16640 1062 16686 1114
rect 16686 1062 16696 1114
rect 16720 1062 16750 1114
rect 16750 1062 16762 1114
rect 16762 1062 16776 1114
rect 16800 1062 16814 1114
rect 16814 1062 16826 1114
rect 16826 1062 16856 1114
rect 16880 1062 16890 1114
rect 16890 1062 16936 1114
rect 16640 1060 16696 1062
rect 16720 1060 16776 1062
rect 16800 1060 16856 1062
rect 16880 1060 16936 1062
rect 24482 1114 24538 1116
rect 24562 1114 24618 1116
rect 24642 1114 24698 1116
rect 24722 1114 24778 1116
rect 24482 1062 24528 1114
rect 24528 1062 24538 1114
rect 24562 1062 24592 1114
rect 24592 1062 24604 1114
rect 24604 1062 24618 1114
rect 24642 1062 24656 1114
rect 24656 1062 24668 1114
rect 24668 1062 24698 1114
rect 24722 1062 24732 1114
rect 24732 1062 24778 1114
rect 24482 1060 24538 1062
rect 24562 1060 24618 1062
rect 24642 1060 24698 1062
rect 24722 1060 24778 1062
rect 32324 1114 32380 1116
rect 32404 1114 32460 1116
rect 32484 1114 32540 1116
rect 32564 1114 32620 1116
rect 32324 1062 32370 1114
rect 32370 1062 32380 1114
rect 32404 1062 32434 1114
rect 32434 1062 32446 1114
rect 32446 1062 32460 1114
rect 32484 1062 32498 1114
rect 32498 1062 32510 1114
rect 32510 1062 32540 1114
rect 32564 1062 32574 1114
rect 32574 1062 32620 1114
rect 32324 1060 32380 1062
rect 32404 1060 32460 1062
rect 32484 1060 32540 1062
rect 32564 1060 32620 1062
<< metal3 >>
rect 2957 21452 3023 21453
rect 4429 21452 4495 21453
rect 2957 21448 3004 21452
rect 3068 21450 3074 21452
rect 2957 21392 2962 21448
rect 2957 21388 3004 21392
rect 3068 21390 3114 21450
rect 4429 21448 4476 21452
rect 4540 21450 4546 21452
rect 4797 21450 4863 21453
rect 5206 21450 5212 21452
rect 4429 21392 4434 21448
rect 3068 21388 3074 21390
rect 4429 21388 4476 21392
rect 4540 21390 4586 21450
rect 4797 21448 5212 21450
rect 4797 21392 4802 21448
rect 4858 21392 5212 21448
rect 4797 21390 5212 21392
rect 4540 21388 4546 21390
rect 2957 21387 3023 21388
rect 4429 21387 4495 21388
rect 4797 21387 4863 21390
rect 5206 21388 5212 21390
rect 5276 21388 5282 21452
rect 5533 21450 5599 21453
rect 5942 21450 5948 21452
rect 5533 21448 5948 21450
rect 5533 21392 5538 21448
rect 5594 21392 5948 21448
rect 5533 21390 5948 21392
rect 5533 21387 5599 21390
rect 5942 21388 5948 21390
rect 6012 21388 6018 21452
rect 6085 21450 6151 21453
rect 8201 21452 8267 21453
rect 9673 21452 9739 21453
rect 6678 21450 6684 21452
rect 6085 21448 6684 21450
rect 6085 21392 6090 21448
rect 6146 21392 6684 21448
rect 6085 21390 6684 21392
rect 6085 21387 6151 21390
rect 6678 21388 6684 21390
rect 6748 21388 6754 21452
rect 8150 21450 8156 21452
rect 8110 21390 8156 21450
rect 8220 21448 8267 21452
rect 8262 21392 8267 21448
rect 8150 21388 8156 21390
rect 8220 21388 8267 21392
rect 9622 21388 9628 21452
rect 9692 21450 9739 21452
rect 9692 21448 9784 21450
rect 9734 21392 9784 21448
rect 9692 21390 9784 21392
rect 9692 21388 9739 21390
rect 11094 21388 11100 21452
rect 11164 21450 11170 21452
rect 11789 21450 11855 21453
rect 11164 21448 11855 21450
rect 11164 21392 11794 21448
rect 11850 21392 11855 21448
rect 11164 21390 11855 21392
rect 11164 21388 11170 21390
rect 8201 21387 8267 21388
rect 9673 21387 9739 21388
rect 11789 21387 11855 21390
rect 13813 21450 13879 21453
rect 14038 21450 14044 21452
rect 13813 21448 14044 21450
rect 13813 21392 13818 21448
rect 13874 21392 14044 21448
rect 13813 21390 14044 21392
rect 13813 21387 13879 21390
rect 14038 21388 14044 21390
rect 14108 21388 14114 21452
rect 14181 21450 14247 21453
rect 14774 21450 14780 21452
rect 14181 21448 14780 21450
rect 14181 21392 14186 21448
rect 14242 21392 14780 21448
rect 14181 21390 14780 21392
rect 14181 21387 14247 21390
rect 14774 21388 14780 21390
rect 14844 21388 14850 21452
rect 15837 21450 15903 21453
rect 16246 21450 16252 21452
rect 15837 21448 16252 21450
rect 15837 21392 15842 21448
rect 15898 21392 16252 21448
rect 15837 21390 16252 21392
rect 15837 21387 15903 21390
rect 16246 21388 16252 21390
rect 16316 21388 16322 21452
rect 28022 21388 28028 21452
rect 28092 21450 28098 21452
rect 28257 21450 28323 21453
rect 28092 21448 28323 21450
rect 28092 21392 28262 21448
rect 28318 21392 28323 21448
rect 28092 21390 28323 21392
rect 28092 21388 28098 21390
rect 28257 21387 28323 21390
rect 28717 21452 28783 21453
rect 29453 21452 29519 21453
rect 28717 21448 28764 21452
rect 28828 21450 28834 21452
rect 28717 21392 28722 21448
rect 28717 21388 28764 21392
rect 28828 21390 28874 21450
rect 29453 21448 29500 21452
rect 29564 21450 29570 21452
rect 29453 21392 29458 21448
rect 28828 21388 28834 21390
rect 29453 21388 29500 21392
rect 29564 21390 29610 21450
rect 29564 21388 29570 21390
rect 30966 21388 30972 21452
rect 31036 21450 31042 21452
rect 31661 21450 31727 21453
rect 31036 21448 31727 21450
rect 31036 21392 31666 21448
rect 31722 21392 31727 21448
rect 31036 21390 31727 21392
rect 31036 21388 31042 21390
rect 28717 21387 28783 21388
rect 29453 21387 29519 21388
rect 31661 21387 31727 21390
rect 10358 21252 10364 21316
rect 10428 21314 10434 21316
rect 11053 21314 11119 21317
rect 10428 21312 11119 21314
rect 10428 21256 11058 21312
rect 11114 21256 11119 21312
rect 10428 21254 11119 21256
rect 10428 21252 10434 21254
rect 11053 21251 11119 21254
rect 11697 21314 11763 21317
rect 11830 21314 11836 21316
rect 11697 21312 11836 21314
rect 11697 21256 11702 21312
rect 11758 21256 11836 21312
rect 11697 21254 11836 21256
rect 11697 21251 11763 21254
rect 11830 21252 11836 21254
rect 11900 21252 11906 21316
rect 12566 21116 12572 21180
rect 12636 21178 12642 21180
rect 13077 21178 13143 21181
rect 12636 21176 13143 21178
rect 12636 21120 13082 21176
rect 13138 21120 13143 21176
rect 12636 21118 13143 21120
rect 12636 21116 12642 21118
rect 13077 21115 13143 21118
rect 27337 21044 27403 21045
rect 27286 21042 27292 21044
rect 27246 20982 27292 21042
rect 27356 21040 27403 21044
rect 27398 20984 27403 21040
rect 27286 20980 27292 20982
rect 27356 20980 27403 20984
rect 27337 20979 27403 20980
rect 8886 20844 8892 20908
rect 8956 20906 8962 20908
rect 9489 20906 9555 20909
rect 8956 20904 9555 20906
rect 8956 20848 9494 20904
rect 9550 20848 9555 20904
rect 8956 20846 9555 20848
rect 8956 20844 8962 20846
rect 9489 20843 9555 20846
rect 16982 20844 16988 20908
rect 17052 20906 17058 20908
rect 17125 20906 17191 20909
rect 17052 20904 17191 20906
rect 17052 20848 17130 20904
rect 17186 20848 17191 20904
rect 17052 20846 17191 20848
rect 17052 20844 17058 20846
rect 17125 20843 17191 20846
rect 8788 20704 9104 20705
rect 8788 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8954 20704
rect 9018 20640 9034 20704
rect 9098 20640 9104 20704
rect 8788 20639 9104 20640
rect 16630 20704 16946 20705
rect 16630 20640 16636 20704
rect 16700 20640 16716 20704
rect 16780 20640 16796 20704
rect 16860 20640 16876 20704
rect 16940 20640 16946 20704
rect 16630 20639 16946 20640
rect 24472 20704 24788 20705
rect 24472 20640 24478 20704
rect 24542 20640 24558 20704
rect 24622 20640 24638 20704
rect 24702 20640 24718 20704
rect 24782 20640 24788 20704
rect 24472 20639 24788 20640
rect 32314 20704 32630 20705
rect 32314 20640 32320 20704
rect 32384 20640 32400 20704
rect 32464 20640 32480 20704
rect 32544 20640 32560 20704
rect 32624 20640 32630 20704
rect 32314 20639 32630 20640
rect 7414 20572 7420 20636
rect 7484 20634 7490 20636
rect 8109 20634 8175 20637
rect 7484 20632 8175 20634
rect 7484 20576 8114 20632
rect 8170 20576 8175 20632
rect 7484 20574 8175 20576
rect 7484 20572 7490 20574
rect 8109 20571 8175 20574
rect 13302 20572 13308 20636
rect 13372 20634 13378 20636
rect 13537 20634 13603 20637
rect 13372 20632 13603 20634
rect 13372 20576 13542 20632
rect 13598 20576 13603 20632
rect 13372 20574 13603 20576
rect 13372 20572 13378 20574
rect 13537 20571 13603 20574
rect 15510 20572 15516 20636
rect 15580 20634 15586 20636
rect 16113 20634 16179 20637
rect 15580 20632 16179 20634
rect 15580 20576 16118 20632
rect 16174 20576 16179 20632
rect 15580 20574 16179 20576
rect 15580 20572 15586 20574
rect 16113 20571 16179 20574
rect 17033 20634 17099 20637
rect 17718 20634 17724 20636
rect 17033 20632 17724 20634
rect 17033 20576 17038 20632
rect 17094 20576 17724 20632
rect 17033 20574 17724 20576
rect 17033 20571 17099 20574
rect 17718 20572 17724 20574
rect 17788 20572 17794 20636
rect 4867 20160 5183 20161
rect 4867 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5113 20160
rect 5177 20096 5183 20160
rect 4867 20095 5183 20096
rect 12709 20160 13025 20161
rect 12709 20096 12715 20160
rect 12779 20096 12795 20160
rect 12859 20096 12875 20160
rect 12939 20096 12955 20160
rect 13019 20096 13025 20160
rect 12709 20095 13025 20096
rect 20551 20160 20867 20161
rect 20551 20096 20557 20160
rect 20621 20096 20637 20160
rect 20701 20096 20717 20160
rect 20781 20096 20797 20160
rect 20861 20096 20867 20160
rect 20551 20095 20867 20096
rect 28393 20160 28709 20161
rect 28393 20096 28399 20160
rect 28463 20096 28479 20160
rect 28543 20096 28559 20160
rect 28623 20096 28639 20160
rect 28703 20096 28709 20160
rect 28393 20095 28709 20096
rect 8788 19616 9104 19617
rect 8788 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8954 19616
rect 9018 19552 9034 19616
rect 9098 19552 9104 19616
rect 8788 19551 9104 19552
rect 16630 19616 16946 19617
rect 16630 19552 16636 19616
rect 16700 19552 16716 19616
rect 16780 19552 16796 19616
rect 16860 19552 16876 19616
rect 16940 19552 16946 19616
rect 16630 19551 16946 19552
rect 24472 19616 24788 19617
rect 24472 19552 24478 19616
rect 24542 19552 24558 19616
rect 24622 19552 24638 19616
rect 24702 19552 24718 19616
rect 24782 19552 24788 19616
rect 24472 19551 24788 19552
rect 32314 19616 32630 19617
rect 32314 19552 32320 19616
rect 32384 19552 32400 19616
rect 32464 19552 32480 19616
rect 32544 19552 32560 19616
rect 32624 19552 32630 19616
rect 32314 19551 32630 19552
rect 1761 19546 1827 19549
rect 2262 19546 2268 19548
rect 1761 19544 2268 19546
rect 1761 19488 1766 19544
rect 1822 19488 2268 19544
rect 1761 19486 2268 19488
rect 1761 19483 1827 19486
rect 2262 19484 2268 19486
rect 2332 19484 2338 19548
rect 18454 19484 18460 19548
rect 18524 19546 18530 19548
rect 18597 19546 18663 19549
rect 18524 19544 18663 19546
rect 18524 19488 18602 19544
rect 18658 19488 18663 19544
rect 18524 19486 18663 19488
rect 18524 19484 18530 19486
rect 18597 19483 18663 19486
rect 13721 19412 13787 19413
rect 13670 19410 13676 19412
rect 13630 19350 13676 19410
rect 13740 19408 13787 19412
rect 13782 19352 13787 19408
rect 13670 19348 13676 19350
rect 13740 19348 13787 19352
rect 13721 19347 13787 19348
rect 19609 19274 19675 19277
rect 22277 19274 22343 19277
rect 19609 19272 22343 19274
rect 19609 19216 19614 19272
rect 19670 19216 22282 19272
rect 22338 19216 22343 19272
rect 19609 19214 22343 19216
rect 19609 19211 19675 19214
rect 22277 19211 22343 19214
rect 4867 19072 5183 19073
rect 4867 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5113 19072
rect 5177 19008 5183 19072
rect 4867 19007 5183 19008
rect 12709 19072 13025 19073
rect 12709 19008 12715 19072
rect 12779 19008 12795 19072
rect 12859 19008 12875 19072
rect 12939 19008 12955 19072
rect 13019 19008 13025 19072
rect 12709 19007 13025 19008
rect 20551 19072 20867 19073
rect 20551 19008 20557 19072
rect 20621 19008 20637 19072
rect 20701 19008 20717 19072
rect 20781 19008 20797 19072
rect 20861 19008 20867 19072
rect 20551 19007 20867 19008
rect 28393 19072 28709 19073
rect 28393 19008 28399 19072
rect 28463 19008 28479 19072
rect 28543 19008 28559 19072
rect 28623 19008 28639 19072
rect 28703 19008 28709 19072
rect 28393 19007 28709 19008
rect 11145 18730 11211 18733
rect 13353 18730 13419 18733
rect 11145 18728 13419 18730
rect 11145 18672 11150 18728
rect 11206 18672 13358 18728
rect 13414 18672 13419 18728
rect 11145 18670 13419 18672
rect 11145 18667 11211 18670
rect 13353 18667 13419 18670
rect 8788 18528 9104 18529
rect 8788 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8954 18528
rect 9018 18464 9034 18528
rect 9098 18464 9104 18528
rect 8788 18463 9104 18464
rect 16630 18528 16946 18529
rect 16630 18464 16636 18528
rect 16700 18464 16716 18528
rect 16780 18464 16796 18528
rect 16860 18464 16876 18528
rect 16940 18464 16946 18528
rect 16630 18463 16946 18464
rect 24472 18528 24788 18529
rect 24472 18464 24478 18528
rect 24542 18464 24558 18528
rect 24622 18464 24638 18528
rect 24702 18464 24718 18528
rect 24782 18464 24788 18528
rect 24472 18463 24788 18464
rect 32314 18528 32630 18529
rect 32314 18464 32320 18528
rect 32384 18464 32400 18528
rect 32464 18464 32480 18528
rect 32544 18464 32560 18528
rect 32624 18464 32630 18528
rect 32314 18463 32630 18464
rect 12341 18186 12407 18189
rect 14181 18186 14247 18189
rect 12341 18184 14247 18186
rect 12341 18128 12346 18184
rect 12402 18128 14186 18184
rect 14242 18128 14247 18184
rect 12341 18126 14247 18128
rect 12341 18123 12407 18126
rect 14181 18123 14247 18126
rect 4867 17984 5183 17985
rect 4867 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5113 17984
rect 5177 17920 5183 17984
rect 4867 17919 5183 17920
rect 12709 17984 13025 17985
rect 12709 17920 12715 17984
rect 12779 17920 12795 17984
rect 12859 17920 12875 17984
rect 12939 17920 12955 17984
rect 13019 17920 13025 17984
rect 12709 17919 13025 17920
rect 20551 17984 20867 17985
rect 20551 17920 20557 17984
rect 20621 17920 20637 17984
rect 20701 17920 20717 17984
rect 20781 17920 20797 17984
rect 20861 17920 20867 17984
rect 20551 17919 20867 17920
rect 28393 17984 28709 17985
rect 28393 17920 28399 17984
rect 28463 17920 28479 17984
rect 28543 17920 28559 17984
rect 28623 17920 28639 17984
rect 28703 17920 28709 17984
rect 28393 17919 28709 17920
rect 1577 17916 1643 17917
rect 1526 17914 1532 17916
rect 1486 17854 1532 17914
rect 1596 17912 1643 17916
rect 1638 17856 1643 17912
rect 1526 17852 1532 17854
rect 1596 17852 1643 17856
rect 1577 17851 1643 17852
rect 3509 17914 3575 17917
rect 3734 17914 3740 17916
rect 3509 17912 3740 17914
rect 3509 17856 3514 17912
rect 3570 17856 3740 17912
rect 3509 17854 3740 17856
rect 3509 17851 3575 17854
rect 3734 17852 3740 17854
rect 3804 17852 3810 17916
rect 15009 17914 15075 17917
rect 14414 17912 15075 17914
rect 14414 17856 15014 17912
rect 15070 17856 15075 17912
rect 14414 17854 15075 17856
rect 11697 17778 11763 17781
rect 14414 17778 14474 17854
rect 15009 17851 15075 17854
rect 15469 17914 15535 17917
rect 16205 17914 16271 17917
rect 15469 17912 16271 17914
rect 15469 17856 15474 17912
rect 15530 17856 16210 17912
rect 16266 17856 16271 17912
rect 15469 17854 16271 17856
rect 15469 17851 15535 17854
rect 16205 17851 16271 17854
rect 21081 17914 21147 17917
rect 25957 17914 26023 17917
rect 21081 17912 26023 17914
rect 21081 17856 21086 17912
rect 21142 17856 25962 17912
rect 26018 17856 26023 17912
rect 21081 17854 26023 17856
rect 21081 17851 21147 17854
rect 25957 17851 26023 17854
rect 31518 17852 31524 17916
rect 31588 17914 31594 17916
rect 31753 17914 31819 17917
rect 31588 17912 31819 17914
rect 31588 17856 31758 17912
rect 31814 17856 31819 17912
rect 31588 17854 31819 17856
rect 31588 17852 31594 17854
rect 31753 17851 31819 17854
rect 11697 17776 14474 17778
rect 11697 17720 11702 17776
rect 11758 17720 14474 17776
rect 11697 17718 14474 17720
rect 14549 17778 14615 17781
rect 25129 17778 25195 17781
rect 14549 17776 25195 17778
rect 14549 17720 14554 17776
rect 14610 17720 25134 17776
rect 25190 17720 25195 17776
rect 14549 17718 25195 17720
rect 11697 17715 11763 17718
rect 14549 17715 14615 17718
rect 25129 17715 25195 17718
rect 7741 17642 7807 17645
rect 26325 17642 26391 17645
rect 7741 17640 26391 17642
rect 7741 17584 7746 17640
rect 7802 17584 26330 17640
rect 26386 17584 26391 17640
rect 7741 17582 26391 17584
rect 7741 17579 7807 17582
rect 26325 17579 26391 17582
rect 13077 17506 13143 17509
rect 15101 17506 15167 17509
rect 13077 17504 15167 17506
rect 13077 17448 13082 17504
rect 13138 17448 15106 17504
rect 15162 17448 15167 17504
rect 13077 17446 15167 17448
rect 13077 17443 13143 17446
rect 15101 17443 15167 17446
rect 8788 17440 9104 17441
rect 8788 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8954 17440
rect 9018 17376 9034 17440
rect 9098 17376 9104 17440
rect 8788 17375 9104 17376
rect 16630 17440 16946 17441
rect 16630 17376 16636 17440
rect 16700 17376 16716 17440
rect 16780 17376 16796 17440
rect 16860 17376 16876 17440
rect 16940 17376 16946 17440
rect 16630 17375 16946 17376
rect 24472 17440 24788 17441
rect 24472 17376 24478 17440
rect 24542 17376 24558 17440
rect 24622 17376 24638 17440
rect 24702 17376 24718 17440
rect 24782 17376 24788 17440
rect 24472 17375 24788 17376
rect 32314 17440 32630 17441
rect 32314 17376 32320 17440
rect 32384 17376 32400 17440
rect 32464 17376 32480 17440
rect 32544 17376 32560 17440
rect 32624 17376 32630 17440
rect 32314 17375 32630 17376
rect 11053 17234 11119 17237
rect 20989 17234 21055 17237
rect 11053 17232 21055 17234
rect 11053 17176 11058 17232
rect 11114 17176 20994 17232
rect 21050 17176 21055 17232
rect 11053 17174 21055 17176
rect 11053 17171 11119 17174
rect 20989 17171 21055 17174
rect 7097 17098 7163 17101
rect 17585 17098 17651 17101
rect 7097 17096 17651 17098
rect 7097 17040 7102 17096
rect 7158 17040 17590 17096
rect 17646 17040 17651 17096
rect 7097 17038 17651 17040
rect 7097 17035 7163 17038
rect 17585 17035 17651 17038
rect 15193 16962 15259 16965
rect 18505 16962 18571 16965
rect 18781 16962 18847 16965
rect 30281 16964 30347 16965
rect 30230 16962 30236 16964
rect 15193 16960 18847 16962
rect 15193 16904 15198 16960
rect 15254 16904 18510 16960
rect 18566 16904 18786 16960
rect 18842 16904 18847 16960
rect 15193 16902 18847 16904
rect 30190 16902 30236 16962
rect 30300 16960 30347 16964
rect 30342 16904 30347 16960
rect 15193 16899 15259 16902
rect 18505 16899 18571 16902
rect 18781 16899 18847 16902
rect 30230 16900 30236 16902
rect 30300 16900 30347 16904
rect 30281 16899 30347 16900
rect 4867 16896 5183 16897
rect 4867 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5113 16896
rect 5177 16832 5183 16896
rect 4867 16831 5183 16832
rect 12709 16896 13025 16897
rect 12709 16832 12715 16896
rect 12779 16832 12795 16896
rect 12859 16832 12875 16896
rect 12939 16832 12955 16896
rect 13019 16832 13025 16896
rect 12709 16831 13025 16832
rect 20551 16896 20867 16897
rect 20551 16832 20557 16896
rect 20621 16832 20637 16896
rect 20701 16832 20717 16896
rect 20781 16832 20797 16896
rect 20861 16832 20867 16896
rect 20551 16831 20867 16832
rect 28393 16896 28709 16897
rect 28393 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28639 16896
rect 28703 16832 28709 16896
rect 28393 16831 28709 16832
rect 10409 16690 10475 16693
rect 16389 16690 16455 16693
rect 10409 16688 16455 16690
rect 10409 16632 10414 16688
rect 10470 16632 16394 16688
rect 16450 16632 16455 16688
rect 10409 16630 16455 16632
rect 10409 16627 10475 16630
rect 16389 16627 16455 16630
rect 14825 16554 14891 16557
rect 19241 16554 19307 16557
rect 14825 16552 19307 16554
rect 14825 16496 14830 16552
rect 14886 16496 19246 16552
rect 19302 16496 19307 16552
rect 14825 16494 19307 16496
rect 14825 16491 14891 16494
rect 19241 16491 19307 16494
rect 21173 16554 21239 16557
rect 23657 16554 23723 16557
rect 21173 16552 23723 16554
rect 21173 16496 21178 16552
rect 21234 16496 23662 16552
rect 23718 16496 23723 16552
rect 21173 16494 23723 16496
rect 21173 16491 21239 16494
rect 23657 16491 23723 16494
rect 18413 16418 18479 16421
rect 20989 16418 21055 16421
rect 18413 16416 21055 16418
rect 18413 16360 18418 16416
rect 18474 16360 20994 16416
rect 21050 16360 21055 16416
rect 18413 16358 21055 16360
rect 18413 16355 18479 16358
rect 20989 16355 21055 16358
rect 8788 16352 9104 16353
rect 8788 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8954 16352
rect 9018 16288 9034 16352
rect 9098 16288 9104 16352
rect 8788 16287 9104 16288
rect 16630 16352 16946 16353
rect 16630 16288 16636 16352
rect 16700 16288 16716 16352
rect 16780 16288 16796 16352
rect 16860 16288 16876 16352
rect 16940 16288 16946 16352
rect 16630 16287 16946 16288
rect 24472 16352 24788 16353
rect 24472 16288 24478 16352
rect 24542 16288 24558 16352
rect 24622 16288 24638 16352
rect 24702 16288 24718 16352
rect 24782 16288 24788 16352
rect 24472 16287 24788 16288
rect 32314 16352 32630 16353
rect 32314 16288 32320 16352
rect 32384 16288 32400 16352
rect 32464 16288 32480 16352
rect 32544 16288 32560 16352
rect 32624 16288 32630 16352
rect 32314 16287 32630 16288
rect 9581 16146 9647 16149
rect 13077 16146 13143 16149
rect 9581 16144 13143 16146
rect 9581 16088 9586 16144
rect 9642 16088 13082 16144
rect 13138 16088 13143 16144
rect 9581 16086 13143 16088
rect 9581 16083 9647 16086
rect 13077 16083 13143 16086
rect 19977 16146 20043 16149
rect 23749 16146 23815 16149
rect 19977 16144 23815 16146
rect 19977 16088 19982 16144
rect 20038 16088 23754 16144
rect 23810 16088 23815 16144
rect 19977 16086 23815 16088
rect 19977 16083 20043 16086
rect 23749 16083 23815 16086
rect 9213 16010 9279 16013
rect 25865 16010 25931 16013
rect 26417 16010 26483 16013
rect 9213 16008 26483 16010
rect 9213 15952 9218 16008
rect 9274 15952 25870 16008
rect 25926 15952 26422 16008
rect 26478 15952 26483 16008
rect 9213 15950 26483 15952
rect 9213 15947 9279 15950
rect 25865 15947 25931 15950
rect 26417 15947 26483 15950
rect 4867 15808 5183 15809
rect 4867 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5113 15808
rect 5177 15744 5183 15808
rect 4867 15743 5183 15744
rect 12709 15808 13025 15809
rect 12709 15744 12715 15808
rect 12779 15744 12795 15808
rect 12859 15744 12875 15808
rect 12939 15744 12955 15808
rect 13019 15744 13025 15808
rect 12709 15743 13025 15744
rect 20551 15808 20867 15809
rect 20551 15744 20557 15808
rect 20621 15744 20637 15808
rect 20701 15744 20717 15808
rect 20781 15744 20797 15808
rect 20861 15744 20867 15808
rect 20551 15743 20867 15744
rect 28393 15808 28709 15809
rect 28393 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28639 15808
rect 28703 15744 28709 15808
rect 28393 15743 28709 15744
rect 19977 15466 20043 15469
rect 21633 15466 21699 15469
rect 19977 15464 21699 15466
rect 19977 15408 19982 15464
rect 20038 15408 21638 15464
rect 21694 15408 21699 15464
rect 19977 15406 21699 15408
rect 19977 15403 20043 15406
rect 21633 15403 21699 15406
rect 23473 15466 23539 15469
rect 25405 15466 25471 15469
rect 23473 15464 25471 15466
rect 23473 15408 23478 15464
rect 23534 15408 25410 15464
rect 25466 15408 25471 15464
rect 23473 15406 25471 15408
rect 23473 15403 23539 15406
rect 25405 15403 25471 15406
rect 21909 15330 21975 15333
rect 23657 15330 23723 15333
rect 21909 15328 23723 15330
rect 21909 15272 21914 15328
rect 21970 15272 23662 15328
rect 23718 15272 23723 15328
rect 21909 15270 23723 15272
rect 21909 15267 21975 15270
rect 23657 15267 23723 15270
rect 8788 15264 9104 15265
rect 8788 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8954 15264
rect 9018 15200 9034 15264
rect 9098 15200 9104 15264
rect 8788 15199 9104 15200
rect 16630 15264 16946 15265
rect 16630 15200 16636 15264
rect 16700 15200 16716 15264
rect 16780 15200 16796 15264
rect 16860 15200 16876 15264
rect 16940 15200 16946 15264
rect 16630 15199 16946 15200
rect 24472 15264 24788 15265
rect 24472 15200 24478 15264
rect 24542 15200 24558 15264
rect 24622 15200 24638 15264
rect 24702 15200 24718 15264
rect 24782 15200 24788 15264
rect 24472 15199 24788 15200
rect 32314 15264 32630 15265
rect 32314 15200 32320 15264
rect 32384 15200 32400 15264
rect 32464 15200 32480 15264
rect 32544 15200 32560 15264
rect 32624 15200 32630 15264
rect 32314 15199 32630 15200
rect 21265 15194 21331 15197
rect 23657 15194 23723 15197
rect 24209 15194 24275 15197
rect 17174 15192 24275 15194
rect 17174 15136 21270 15192
rect 21326 15136 23662 15192
rect 23718 15136 24214 15192
rect 24270 15136 24275 15192
rect 17174 15134 24275 15136
rect 13721 15058 13787 15061
rect 17174 15058 17234 15134
rect 21265 15131 21331 15134
rect 23657 15131 23723 15134
rect 24209 15131 24275 15134
rect 13721 15056 17234 15058
rect 13721 15000 13726 15056
rect 13782 15000 17234 15056
rect 13721 14998 17234 15000
rect 13721 14995 13787 14998
rect 8661 14922 8727 14925
rect 22185 14922 22251 14925
rect 8661 14920 22251 14922
rect 8661 14864 8666 14920
rect 8722 14864 22190 14920
rect 22246 14864 22251 14920
rect 8661 14862 22251 14864
rect 8661 14859 8727 14862
rect 22185 14859 22251 14862
rect 4867 14720 5183 14721
rect 4867 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5113 14720
rect 5177 14656 5183 14720
rect 4867 14655 5183 14656
rect 12709 14720 13025 14721
rect 12709 14656 12715 14720
rect 12779 14656 12795 14720
rect 12859 14656 12875 14720
rect 12939 14656 12955 14720
rect 13019 14656 13025 14720
rect 12709 14655 13025 14656
rect 20551 14720 20867 14721
rect 20551 14656 20557 14720
rect 20621 14656 20637 14720
rect 20701 14656 20717 14720
rect 20781 14656 20797 14720
rect 20861 14656 20867 14720
rect 20551 14655 20867 14656
rect 28393 14720 28709 14721
rect 28393 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28639 14720
rect 28703 14656 28709 14720
rect 28393 14655 28709 14656
rect 12709 14514 12775 14517
rect 14365 14514 14431 14517
rect 12709 14512 14431 14514
rect 12709 14456 12714 14512
rect 12770 14456 14370 14512
rect 14426 14456 14431 14512
rect 12709 14454 14431 14456
rect 12709 14451 12775 14454
rect 14365 14451 14431 14454
rect 26233 14514 26299 14517
rect 28717 14514 28783 14517
rect 26233 14512 28783 14514
rect 26233 14456 26238 14512
rect 26294 14456 28722 14512
rect 28778 14456 28783 14512
rect 26233 14454 28783 14456
rect 26233 14451 26299 14454
rect 28717 14451 28783 14454
rect 25957 14378 26023 14381
rect 28809 14378 28875 14381
rect 25957 14376 28875 14378
rect 25957 14320 25962 14376
rect 26018 14320 28814 14376
rect 28870 14320 28875 14376
rect 25957 14318 28875 14320
rect 25957 14315 26023 14318
rect 28809 14315 28875 14318
rect 8788 14176 9104 14177
rect 8788 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8954 14176
rect 9018 14112 9034 14176
rect 9098 14112 9104 14176
rect 8788 14111 9104 14112
rect 16630 14176 16946 14177
rect 16630 14112 16636 14176
rect 16700 14112 16716 14176
rect 16780 14112 16796 14176
rect 16860 14112 16876 14176
rect 16940 14112 16946 14176
rect 16630 14111 16946 14112
rect 24472 14176 24788 14177
rect 24472 14112 24478 14176
rect 24542 14112 24558 14176
rect 24622 14112 24638 14176
rect 24702 14112 24718 14176
rect 24782 14112 24788 14176
rect 24472 14111 24788 14112
rect 32314 14176 32630 14177
rect 32314 14112 32320 14176
rect 32384 14112 32400 14176
rect 32464 14112 32480 14176
rect 32544 14112 32560 14176
rect 32624 14112 32630 14176
rect 32314 14111 32630 14112
rect 13077 13970 13143 13973
rect 18413 13970 18479 13973
rect 13077 13968 18479 13970
rect 13077 13912 13082 13968
rect 13138 13912 18418 13968
rect 18474 13912 18479 13968
rect 13077 13910 18479 13912
rect 13077 13907 13143 13910
rect 18413 13907 18479 13910
rect 20161 13834 20227 13837
rect 24209 13834 24275 13837
rect 20161 13832 24275 13834
rect 20161 13776 20166 13832
rect 20222 13776 24214 13832
rect 24270 13776 24275 13832
rect 20161 13774 24275 13776
rect 20161 13771 20227 13774
rect 24209 13771 24275 13774
rect 4867 13632 5183 13633
rect 4867 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5113 13632
rect 5177 13568 5183 13632
rect 4867 13567 5183 13568
rect 12709 13632 13025 13633
rect 12709 13568 12715 13632
rect 12779 13568 12795 13632
rect 12859 13568 12875 13632
rect 12939 13568 12955 13632
rect 13019 13568 13025 13632
rect 12709 13567 13025 13568
rect 20551 13632 20867 13633
rect 20551 13568 20557 13632
rect 20621 13568 20637 13632
rect 20701 13568 20717 13632
rect 20781 13568 20797 13632
rect 20861 13568 20867 13632
rect 20551 13567 20867 13568
rect 28393 13632 28709 13633
rect 28393 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28639 13632
rect 28703 13568 28709 13632
rect 28393 13567 28709 13568
rect 11513 13426 11579 13429
rect 22001 13426 22067 13429
rect 11513 13424 22067 13426
rect 11513 13368 11518 13424
rect 11574 13368 22006 13424
rect 22062 13368 22067 13424
rect 11513 13366 22067 13368
rect 11513 13363 11579 13366
rect 22001 13363 22067 13366
rect 14641 13290 14707 13293
rect 24669 13290 24735 13293
rect 14641 13288 24735 13290
rect 14641 13232 14646 13288
rect 14702 13232 24674 13288
rect 24730 13232 24735 13288
rect 14641 13230 24735 13232
rect 14641 13227 14707 13230
rect 24669 13227 24735 13230
rect 8788 13088 9104 13089
rect 8788 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8954 13088
rect 9018 13024 9034 13088
rect 9098 13024 9104 13088
rect 8788 13023 9104 13024
rect 16630 13088 16946 13089
rect 16630 13024 16636 13088
rect 16700 13024 16716 13088
rect 16780 13024 16796 13088
rect 16860 13024 16876 13088
rect 16940 13024 16946 13088
rect 16630 13023 16946 13024
rect 24472 13088 24788 13089
rect 24472 13024 24478 13088
rect 24542 13024 24558 13088
rect 24622 13024 24638 13088
rect 24702 13024 24718 13088
rect 24782 13024 24788 13088
rect 24472 13023 24788 13024
rect 32314 13088 32630 13089
rect 32314 13024 32320 13088
rect 32384 13024 32400 13088
rect 32464 13024 32480 13088
rect 32544 13024 32560 13088
rect 32624 13024 32630 13088
rect 32314 13023 32630 13024
rect 13169 13018 13235 13021
rect 14733 13018 14799 13021
rect 15561 13018 15627 13021
rect 13169 13016 15627 13018
rect 13169 12960 13174 13016
rect 13230 12960 14738 13016
rect 14794 12960 15566 13016
rect 15622 12960 15627 13016
rect 13169 12958 15627 12960
rect 13169 12955 13235 12958
rect 14733 12955 14799 12958
rect 15561 12955 15627 12958
rect 4867 12544 5183 12545
rect 4867 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5113 12544
rect 5177 12480 5183 12544
rect 4867 12479 5183 12480
rect 12709 12544 13025 12545
rect 12709 12480 12715 12544
rect 12779 12480 12795 12544
rect 12859 12480 12875 12544
rect 12939 12480 12955 12544
rect 13019 12480 13025 12544
rect 12709 12479 13025 12480
rect 20551 12544 20867 12545
rect 20551 12480 20557 12544
rect 20621 12480 20637 12544
rect 20701 12480 20717 12544
rect 20781 12480 20797 12544
rect 20861 12480 20867 12544
rect 20551 12479 20867 12480
rect 28393 12544 28709 12545
rect 28393 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28639 12544
rect 28703 12480 28709 12544
rect 28393 12479 28709 12480
rect 13670 12276 13676 12340
rect 13740 12338 13746 12340
rect 14273 12338 14339 12341
rect 13740 12336 14339 12338
rect 13740 12280 14278 12336
rect 14334 12280 14339 12336
rect 13740 12278 14339 12280
rect 13740 12276 13746 12278
rect 14273 12275 14339 12278
rect 8788 12000 9104 12001
rect 8788 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8954 12000
rect 9018 11936 9034 12000
rect 9098 11936 9104 12000
rect 8788 11935 9104 11936
rect 16630 12000 16946 12001
rect 16630 11936 16636 12000
rect 16700 11936 16716 12000
rect 16780 11936 16796 12000
rect 16860 11936 16876 12000
rect 16940 11936 16946 12000
rect 16630 11935 16946 11936
rect 24472 12000 24788 12001
rect 24472 11936 24478 12000
rect 24542 11936 24558 12000
rect 24622 11936 24638 12000
rect 24702 11936 24718 12000
rect 24782 11936 24788 12000
rect 24472 11935 24788 11936
rect 32314 12000 32630 12001
rect 32314 11936 32320 12000
rect 32384 11936 32400 12000
rect 32464 11936 32480 12000
rect 32544 11936 32560 12000
rect 32624 11936 32630 12000
rect 32314 11935 32630 11936
rect 14457 11794 14523 11797
rect 18781 11794 18847 11797
rect 14457 11792 18847 11794
rect 14457 11736 14462 11792
rect 14518 11736 18786 11792
rect 18842 11736 18847 11792
rect 14457 11734 18847 11736
rect 14457 11731 14523 11734
rect 18781 11731 18847 11734
rect 4867 11456 5183 11457
rect 4867 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5113 11456
rect 5177 11392 5183 11456
rect 4867 11391 5183 11392
rect 12709 11456 13025 11457
rect 12709 11392 12715 11456
rect 12779 11392 12795 11456
rect 12859 11392 12875 11456
rect 12939 11392 12955 11456
rect 13019 11392 13025 11456
rect 12709 11391 13025 11392
rect 20551 11456 20867 11457
rect 20551 11392 20557 11456
rect 20621 11392 20637 11456
rect 20701 11392 20717 11456
rect 20781 11392 20797 11456
rect 20861 11392 20867 11456
rect 20551 11391 20867 11392
rect 28393 11456 28709 11457
rect 28393 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28639 11456
rect 28703 11392 28709 11456
rect 28393 11391 28709 11392
rect 13629 11114 13695 11117
rect 16941 11114 17007 11117
rect 13629 11112 17007 11114
rect 13629 11056 13634 11112
rect 13690 11056 16946 11112
rect 17002 11056 17007 11112
rect 13629 11054 17007 11056
rect 13629 11051 13695 11054
rect 16941 11051 17007 11054
rect 8788 10912 9104 10913
rect 8788 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8954 10912
rect 9018 10848 9034 10912
rect 9098 10848 9104 10912
rect 8788 10847 9104 10848
rect 16630 10912 16946 10913
rect 16630 10848 16636 10912
rect 16700 10848 16716 10912
rect 16780 10848 16796 10912
rect 16860 10848 16876 10912
rect 16940 10848 16946 10912
rect 16630 10847 16946 10848
rect 24472 10912 24788 10913
rect 24472 10848 24478 10912
rect 24542 10848 24558 10912
rect 24622 10848 24638 10912
rect 24702 10848 24718 10912
rect 24782 10848 24788 10912
rect 24472 10847 24788 10848
rect 32314 10912 32630 10913
rect 32314 10848 32320 10912
rect 32384 10848 32400 10912
rect 32464 10848 32480 10912
rect 32544 10848 32560 10912
rect 32624 10848 32630 10912
rect 32314 10847 32630 10848
rect 4867 10368 5183 10369
rect 4867 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5113 10368
rect 5177 10304 5183 10368
rect 4867 10303 5183 10304
rect 12709 10368 13025 10369
rect 12709 10304 12715 10368
rect 12779 10304 12795 10368
rect 12859 10304 12875 10368
rect 12939 10304 12955 10368
rect 13019 10304 13025 10368
rect 12709 10303 13025 10304
rect 20551 10368 20867 10369
rect 20551 10304 20557 10368
rect 20621 10304 20637 10368
rect 20701 10304 20717 10368
rect 20781 10304 20797 10368
rect 20861 10304 20867 10368
rect 20551 10303 20867 10304
rect 28393 10368 28709 10369
rect 28393 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28639 10368
rect 28703 10304 28709 10368
rect 28393 10303 28709 10304
rect 8788 9824 9104 9825
rect 8788 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8954 9824
rect 9018 9760 9034 9824
rect 9098 9760 9104 9824
rect 8788 9759 9104 9760
rect 16630 9824 16946 9825
rect 16630 9760 16636 9824
rect 16700 9760 16716 9824
rect 16780 9760 16796 9824
rect 16860 9760 16876 9824
rect 16940 9760 16946 9824
rect 16630 9759 16946 9760
rect 24472 9824 24788 9825
rect 24472 9760 24478 9824
rect 24542 9760 24558 9824
rect 24622 9760 24638 9824
rect 24702 9760 24718 9824
rect 24782 9760 24788 9824
rect 24472 9759 24788 9760
rect 32314 9824 32630 9825
rect 32314 9760 32320 9824
rect 32384 9760 32400 9824
rect 32464 9760 32480 9824
rect 32544 9760 32560 9824
rect 32624 9760 32630 9824
rect 32314 9759 32630 9760
rect 9673 9618 9739 9621
rect 10409 9618 10475 9621
rect 11421 9618 11487 9621
rect 13537 9618 13603 9621
rect 9673 9616 13603 9618
rect 9673 9560 9678 9616
rect 9734 9560 10414 9616
rect 10470 9560 11426 9616
rect 11482 9560 13542 9616
rect 13598 9560 13603 9616
rect 9673 9558 13603 9560
rect 9673 9555 9739 9558
rect 10409 9555 10475 9558
rect 11421 9555 11487 9558
rect 13537 9555 13603 9558
rect 4867 9280 5183 9281
rect 4867 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5113 9280
rect 5177 9216 5183 9280
rect 4867 9215 5183 9216
rect 12709 9280 13025 9281
rect 12709 9216 12715 9280
rect 12779 9216 12795 9280
rect 12859 9216 12875 9280
rect 12939 9216 12955 9280
rect 13019 9216 13025 9280
rect 12709 9215 13025 9216
rect 20551 9280 20867 9281
rect 20551 9216 20557 9280
rect 20621 9216 20637 9280
rect 20701 9216 20717 9280
rect 20781 9216 20797 9280
rect 20861 9216 20867 9280
rect 20551 9215 20867 9216
rect 28393 9280 28709 9281
rect 28393 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28639 9280
rect 28703 9216 28709 9280
rect 28393 9215 28709 9216
rect 20713 9074 20779 9077
rect 25405 9074 25471 9077
rect 26969 9074 27035 9077
rect 20713 9072 27035 9074
rect 20713 9016 20718 9072
rect 20774 9016 25410 9072
rect 25466 9016 26974 9072
rect 27030 9016 27035 9072
rect 20713 9014 27035 9016
rect 20713 9011 20779 9014
rect 25405 9011 25471 9014
rect 26969 9011 27035 9014
rect 5901 8938 5967 8941
rect 13629 8938 13695 8941
rect 5901 8936 13695 8938
rect 5901 8880 5906 8936
rect 5962 8880 13634 8936
rect 13690 8880 13695 8936
rect 5901 8878 13695 8880
rect 5901 8875 5967 8878
rect 13629 8875 13695 8878
rect 8788 8736 9104 8737
rect 8788 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8954 8736
rect 9018 8672 9034 8736
rect 9098 8672 9104 8736
rect 8788 8671 9104 8672
rect 16630 8736 16946 8737
rect 16630 8672 16636 8736
rect 16700 8672 16716 8736
rect 16780 8672 16796 8736
rect 16860 8672 16876 8736
rect 16940 8672 16946 8736
rect 16630 8671 16946 8672
rect 24472 8736 24788 8737
rect 24472 8672 24478 8736
rect 24542 8672 24558 8736
rect 24622 8672 24638 8736
rect 24702 8672 24718 8736
rect 24782 8672 24788 8736
rect 24472 8671 24788 8672
rect 32314 8736 32630 8737
rect 32314 8672 32320 8736
rect 32384 8672 32400 8736
rect 32464 8672 32480 8736
rect 32544 8672 32560 8736
rect 32624 8672 32630 8736
rect 32314 8671 32630 8672
rect 10133 8530 10199 8533
rect 14181 8530 14247 8533
rect 10133 8528 14247 8530
rect 10133 8472 10138 8528
rect 10194 8472 14186 8528
rect 14242 8472 14247 8528
rect 10133 8470 14247 8472
rect 10133 8467 10199 8470
rect 14181 8467 14247 8470
rect 4867 8192 5183 8193
rect 4867 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5113 8192
rect 5177 8128 5183 8192
rect 4867 8127 5183 8128
rect 12709 8192 13025 8193
rect 12709 8128 12715 8192
rect 12779 8128 12795 8192
rect 12859 8128 12875 8192
rect 12939 8128 12955 8192
rect 13019 8128 13025 8192
rect 12709 8127 13025 8128
rect 20551 8192 20867 8193
rect 20551 8128 20557 8192
rect 20621 8128 20637 8192
rect 20701 8128 20717 8192
rect 20781 8128 20797 8192
rect 20861 8128 20867 8192
rect 20551 8127 20867 8128
rect 28393 8192 28709 8193
rect 28393 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28639 8192
rect 28703 8128 28709 8192
rect 28393 8127 28709 8128
rect 8788 7648 9104 7649
rect 8788 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8954 7648
rect 9018 7584 9034 7648
rect 9098 7584 9104 7648
rect 8788 7583 9104 7584
rect 16630 7648 16946 7649
rect 16630 7584 16636 7648
rect 16700 7584 16716 7648
rect 16780 7584 16796 7648
rect 16860 7584 16876 7648
rect 16940 7584 16946 7648
rect 16630 7583 16946 7584
rect 24472 7648 24788 7649
rect 24472 7584 24478 7648
rect 24542 7584 24558 7648
rect 24622 7584 24638 7648
rect 24702 7584 24718 7648
rect 24782 7584 24788 7648
rect 24472 7583 24788 7584
rect 32314 7648 32630 7649
rect 32314 7584 32320 7648
rect 32384 7584 32400 7648
rect 32464 7584 32480 7648
rect 32544 7584 32560 7648
rect 32624 7584 32630 7648
rect 32314 7583 32630 7584
rect 4867 7104 5183 7105
rect 4867 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5113 7104
rect 5177 7040 5183 7104
rect 4867 7039 5183 7040
rect 12709 7104 13025 7105
rect 12709 7040 12715 7104
rect 12779 7040 12795 7104
rect 12859 7040 12875 7104
rect 12939 7040 12955 7104
rect 13019 7040 13025 7104
rect 12709 7039 13025 7040
rect 20551 7104 20867 7105
rect 20551 7040 20557 7104
rect 20621 7040 20637 7104
rect 20701 7040 20717 7104
rect 20781 7040 20797 7104
rect 20861 7040 20867 7104
rect 20551 7039 20867 7040
rect 28393 7104 28709 7105
rect 28393 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28639 7104
rect 28703 7040 28709 7104
rect 28393 7039 28709 7040
rect 8788 6560 9104 6561
rect 8788 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8954 6560
rect 9018 6496 9034 6560
rect 9098 6496 9104 6560
rect 8788 6495 9104 6496
rect 16630 6560 16946 6561
rect 16630 6496 16636 6560
rect 16700 6496 16716 6560
rect 16780 6496 16796 6560
rect 16860 6496 16876 6560
rect 16940 6496 16946 6560
rect 16630 6495 16946 6496
rect 24472 6560 24788 6561
rect 24472 6496 24478 6560
rect 24542 6496 24558 6560
rect 24622 6496 24638 6560
rect 24702 6496 24718 6560
rect 24782 6496 24788 6560
rect 24472 6495 24788 6496
rect 32314 6560 32630 6561
rect 32314 6496 32320 6560
rect 32384 6496 32400 6560
rect 32464 6496 32480 6560
rect 32544 6496 32560 6560
rect 32624 6496 32630 6560
rect 32314 6495 32630 6496
rect 4867 6016 5183 6017
rect 4867 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5113 6016
rect 5177 5952 5183 6016
rect 4867 5951 5183 5952
rect 12709 6016 13025 6017
rect 12709 5952 12715 6016
rect 12779 5952 12795 6016
rect 12859 5952 12875 6016
rect 12939 5952 12955 6016
rect 13019 5952 13025 6016
rect 12709 5951 13025 5952
rect 20551 6016 20867 6017
rect 20551 5952 20557 6016
rect 20621 5952 20637 6016
rect 20701 5952 20717 6016
rect 20781 5952 20797 6016
rect 20861 5952 20867 6016
rect 20551 5951 20867 5952
rect 28393 6016 28709 6017
rect 28393 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28639 6016
rect 28703 5952 28709 6016
rect 28393 5951 28709 5952
rect 8788 5472 9104 5473
rect 8788 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8954 5472
rect 9018 5408 9034 5472
rect 9098 5408 9104 5472
rect 8788 5407 9104 5408
rect 16630 5472 16946 5473
rect 16630 5408 16636 5472
rect 16700 5408 16716 5472
rect 16780 5408 16796 5472
rect 16860 5408 16876 5472
rect 16940 5408 16946 5472
rect 16630 5407 16946 5408
rect 24472 5472 24788 5473
rect 24472 5408 24478 5472
rect 24542 5408 24558 5472
rect 24622 5408 24638 5472
rect 24702 5408 24718 5472
rect 24782 5408 24788 5472
rect 24472 5407 24788 5408
rect 32314 5472 32630 5473
rect 32314 5408 32320 5472
rect 32384 5408 32400 5472
rect 32464 5408 32480 5472
rect 32544 5408 32560 5472
rect 32624 5408 32630 5472
rect 32314 5407 32630 5408
rect 4867 4928 5183 4929
rect 4867 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5113 4928
rect 5177 4864 5183 4928
rect 4867 4863 5183 4864
rect 12709 4928 13025 4929
rect 12709 4864 12715 4928
rect 12779 4864 12795 4928
rect 12859 4864 12875 4928
rect 12939 4864 12955 4928
rect 13019 4864 13025 4928
rect 12709 4863 13025 4864
rect 20551 4928 20867 4929
rect 20551 4864 20557 4928
rect 20621 4864 20637 4928
rect 20701 4864 20717 4928
rect 20781 4864 20797 4928
rect 20861 4864 20867 4928
rect 20551 4863 20867 4864
rect 28393 4928 28709 4929
rect 28393 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28639 4928
rect 28703 4864 28709 4928
rect 28393 4863 28709 4864
rect 8788 4384 9104 4385
rect 8788 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8954 4384
rect 9018 4320 9034 4384
rect 9098 4320 9104 4384
rect 8788 4319 9104 4320
rect 16630 4384 16946 4385
rect 16630 4320 16636 4384
rect 16700 4320 16716 4384
rect 16780 4320 16796 4384
rect 16860 4320 16876 4384
rect 16940 4320 16946 4384
rect 16630 4319 16946 4320
rect 24472 4384 24788 4385
rect 24472 4320 24478 4384
rect 24542 4320 24558 4384
rect 24622 4320 24638 4384
rect 24702 4320 24718 4384
rect 24782 4320 24788 4384
rect 24472 4319 24788 4320
rect 32314 4384 32630 4385
rect 32314 4320 32320 4384
rect 32384 4320 32400 4384
rect 32464 4320 32480 4384
rect 32544 4320 32560 4384
rect 32624 4320 32630 4384
rect 32314 4319 32630 4320
rect 4867 3840 5183 3841
rect 4867 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5113 3840
rect 5177 3776 5183 3840
rect 4867 3775 5183 3776
rect 12709 3840 13025 3841
rect 12709 3776 12715 3840
rect 12779 3776 12795 3840
rect 12859 3776 12875 3840
rect 12939 3776 12955 3840
rect 13019 3776 13025 3840
rect 12709 3775 13025 3776
rect 20551 3840 20867 3841
rect 20551 3776 20557 3840
rect 20621 3776 20637 3840
rect 20701 3776 20717 3840
rect 20781 3776 20797 3840
rect 20861 3776 20867 3840
rect 20551 3775 20867 3776
rect 28393 3840 28709 3841
rect 28393 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28639 3840
rect 28703 3776 28709 3840
rect 28393 3775 28709 3776
rect 8788 3296 9104 3297
rect 8788 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8954 3296
rect 9018 3232 9034 3296
rect 9098 3232 9104 3296
rect 8788 3231 9104 3232
rect 16630 3296 16946 3297
rect 16630 3232 16636 3296
rect 16700 3232 16716 3296
rect 16780 3232 16796 3296
rect 16860 3232 16876 3296
rect 16940 3232 16946 3296
rect 16630 3231 16946 3232
rect 24472 3296 24788 3297
rect 24472 3232 24478 3296
rect 24542 3232 24558 3296
rect 24622 3232 24638 3296
rect 24702 3232 24718 3296
rect 24782 3232 24788 3296
rect 24472 3231 24788 3232
rect 32314 3296 32630 3297
rect 32314 3232 32320 3296
rect 32384 3232 32400 3296
rect 32464 3232 32480 3296
rect 32544 3232 32560 3296
rect 32624 3232 32630 3296
rect 32314 3231 32630 3232
rect 4867 2752 5183 2753
rect 4867 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5113 2752
rect 5177 2688 5183 2752
rect 4867 2687 5183 2688
rect 12709 2752 13025 2753
rect 12709 2688 12715 2752
rect 12779 2688 12795 2752
rect 12859 2688 12875 2752
rect 12939 2688 12955 2752
rect 13019 2688 13025 2752
rect 12709 2687 13025 2688
rect 20551 2752 20867 2753
rect 20551 2688 20557 2752
rect 20621 2688 20637 2752
rect 20701 2688 20717 2752
rect 20781 2688 20797 2752
rect 20861 2688 20867 2752
rect 20551 2687 20867 2688
rect 28393 2752 28709 2753
rect 28393 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28639 2752
rect 28703 2688 28709 2752
rect 28393 2687 28709 2688
rect 8788 2208 9104 2209
rect 8788 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8954 2208
rect 9018 2144 9034 2208
rect 9098 2144 9104 2208
rect 8788 2143 9104 2144
rect 16630 2208 16946 2209
rect 16630 2144 16636 2208
rect 16700 2144 16716 2208
rect 16780 2144 16796 2208
rect 16860 2144 16876 2208
rect 16940 2144 16946 2208
rect 16630 2143 16946 2144
rect 24472 2208 24788 2209
rect 24472 2144 24478 2208
rect 24542 2144 24558 2208
rect 24622 2144 24638 2208
rect 24702 2144 24718 2208
rect 24782 2144 24788 2208
rect 24472 2143 24788 2144
rect 32314 2208 32630 2209
rect 32314 2144 32320 2208
rect 32384 2144 32400 2208
rect 32464 2144 32480 2208
rect 32544 2144 32560 2208
rect 32624 2144 32630 2208
rect 32314 2143 32630 2144
rect 4867 1664 5183 1665
rect 4867 1600 4873 1664
rect 4937 1600 4953 1664
rect 5017 1600 5033 1664
rect 5097 1600 5113 1664
rect 5177 1600 5183 1664
rect 4867 1599 5183 1600
rect 12709 1664 13025 1665
rect 12709 1600 12715 1664
rect 12779 1600 12795 1664
rect 12859 1600 12875 1664
rect 12939 1600 12955 1664
rect 13019 1600 13025 1664
rect 12709 1599 13025 1600
rect 20551 1664 20867 1665
rect 20551 1600 20557 1664
rect 20621 1600 20637 1664
rect 20701 1600 20717 1664
rect 20781 1600 20797 1664
rect 20861 1600 20867 1664
rect 20551 1599 20867 1600
rect 28393 1664 28709 1665
rect 28393 1600 28399 1664
rect 28463 1600 28479 1664
rect 28543 1600 28559 1664
rect 28623 1600 28639 1664
rect 28703 1600 28709 1664
rect 28393 1599 28709 1600
rect 8788 1120 9104 1121
rect 8788 1056 8794 1120
rect 8858 1056 8874 1120
rect 8938 1056 8954 1120
rect 9018 1056 9034 1120
rect 9098 1056 9104 1120
rect 8788 1055 9104 1056
rect 16630 1120 16946 1121
rect 16630 1056 16636 1120
rect 16700 1056 16716 1120
rect 16780 1056 16796 1120
rect 16860 1056 16876 1120
rect 16940 1056 16946 1120
rect 16630 1055 16946 1056
rect 24472 1120 24788 1121
rect 24472 1056 24478 1120
rect 24542 1056 24558 1120
rect 24622 1056 24638 1120
rect 24702 1056 24718 1120
rect 24782 1056 24788 1120
rect 24472 1055 24788 1056
rect 32314 1120 32630 1121
rect 32314 1056 32320 1120
rect 32384 1056 32400 1120
rect 32464 1056 32480 1120
rect 32544 1056 32560 1120
rect 32624 1056 32630 1120
rect 32314 1055 32630 1056
<< via3 >>
rect 3004 21448 3068 21452
rect 3004 21392 3018 21448
rect 3018 21392 3068 21448
rect 3004 21388 3068 21392
rect 4476 21448 4540 21452
rect 4476 21392 4490 21448
rect 4490 21392 4540 21448
rect 4476 21388 4540 21392
rect 5212 21388 5276 21452
rect 5948 21388 6012 21452
rect 6684 21388 6748 21452
rect 8156 21448 8220 21452
rect 8156 21392 8206 21448
rect 8206 21392 8220 21448
rect 8156 21388 8220 21392
rect 9628 21448 9692 21452
rect 9628 21392 9678 21448
rect 9678 21392 9692 21448
rect 9628 21388 9692 21392
rect 11100 21388 11164 21452
rect 14044 21388 14108 21452
rect 14780 21388 14844 21452
rect 16252 21388 16316 21452
rect 28028 21388 28092 21452
rect 28764 21448 28828 21452
rect 28764 21392 28778 21448
rect 28778 21392 28828 21448
rect 28764 21388 28828 21392
rect 29500 21448 29564 21452
rect 29500 21392 29514 21448
rect 29514 21392 29564 21448
rect 29500 21388 29564 21392
rect 30972 21388 31036 21452
rect 10364 21252 10428 21316
rect 11836 21252 11900 21316
rect 12572 21116 12636 21180
rect 27292 21040 27356 21044
rect 27292 20984 27342 21040
rect 27342 20984 27356 21040
rect 27292 20980 27356 20984
rect 8892 20844 8956 20908
rect 16988 20844 17052 20908
rect 8794 20700 8858 20704
rect 8794 20644 8798 20700
rect 8798 20644 8854 20700
rect 8854 20644 8858 20700
rect 8794 20640 8858 20644
rect 8874 20700 8938 20704
rect 8874 20644 8878 20700
rect 8878 20644 8934 20700
rect 8934 20644 8938 20700
rect 8874 20640 8938 20644
rect 8954 20700 9018 20704
rect 8954 20644 8958 20700
rect 8958 20644 9014 20700
rect 9014 20644 9018 20700
rect 8954 20640 9018 20644
rect 9034 20700 9098 20704
rect 9034 20644 9038 20700
rect 9038 20644 9094 20700
rect 9094 20644 9098 20700
rect 9034 20640 9098 20644
rect 16636 20700 16700 20704
rect 16636 20644 16640 20700
rect 16640 20644 16696 20700
rect 16696 20644 16700 20700
rect 16636 20640 16700 20644
rect 16716 20700 16780 20704
rect 16716 20644 16720 20700
rect 16720 20644 16776 20700
rect 16776 20644 16780 20700
rect 16716 20640 16780 20644
rect 16796 20700 16860 20704
rect 16796 20644 16800 20700
rect 16800 20644 16856 20700
rect 16856 20644 16860 20700
rect 16796 20640 16860 20644
rect 16876 20700 16940 20704
rect 16876 20644 16880 20700
rect 16880 20644 16936 20700
rect 16936 20644 16940 20700
rect 16876 20640 16940 20644
rect 24478 20700 24542 20704
rect 24478 20644 24482 20700
rect 24482 20644 24538 20700
rect 24538 20644 24542 20700
rect 24478 20640 24542 20644
rect 24558 20700 24622 20704
rect 24558 20644 24562 20700
rect 24562 20644 24618 20700
rect 24618 20644 24622 20700
rect 24558 20640 24622 20644
rect 24638 20700 24702 20704
rect 24638 20644 24642 20700
rect 24642 20644 24698 20700
rect 24698 20644 24702 20700
rect 24638 20640 24702 20644
rect 24718 20700 24782 20704
rect 24718 20644 24722 20700
rect 24722 20644 24778 20700
rect 24778 20644 24782 20700
rect 24718 20640 24782 20644
rect 32320 20700 32384 20704
rect 32320 20644 32324 20700
rect 32324 20644 32380 20700
rect 32380 20644 32384 20700
rect 32320 20640 32384 20644
rect 32400 20700 32464 20704
rect 32400 20644 32404 20700
rect 32404 20644 32460 20700
rect 32460 20644 32464 20700
rect 32400 20640 32464 20644
rect 32480 20700 32544 20704
rect 32480 20644 32484 20700
rect 32484 20644 32540 20700
rect 32540 20644 32544 20700
rect 32480 20640 32544 20644
rect 32560 20700 32624 20704
rect 32560 20644 32564 20700
rect 32564 20644 32620 20700
rect 32620 20644 32624 20700
rect 32560 20640 32624 20644
rect 7420 20572 7484 20636
rect 13308 20572 13372 20636
rect 15516 20572 15580 20636
rect 17724 20572 17788 20636
rect 4873 20156 4937 20160
rect 4873 20100 4877 20156
rect 4877 20100 4933 20156
rect 4933 20100 4937 20156
rect 4873 20096 4937 20100
rect 4953 20156 5017 20160
rect 4953 20100 4957 20156
rect 4957 20100 5013 20156
rect 5013 20100 5017 20156
rect 4953 20096 5017 20100
rect 5033 20156 5097 20160
rect 5033 20100 5037 20156
rect 5037 20100 5093 20156
rect 5093 20100 5097 20156
rect 5033 20096 5097 20100
rect 5113 20156 5177 20160
rect 5113 20100 5117 20156
rect 5117 20100 5173 20156
rect 5173 20100 5177 20156
rect 5113 20096 5177 20100
rect 12715 20156 12779 20160
rect 12715 20100 12719 20156
rect 12719 20100 12775 20156
rect 12775 20100 12779 20156
rect 12715 20096 12779 20100
rect 12795 20156 12859 20160
rect 12795 20100 12799 20156
rect 12799 20100 12855 20156
rect 12855 20100 12859 20156
rect 12795 20096 12859 20100
rect 12875 20156 12939 20160
rect 12875 20100 12879 20156
rect 12879 20100 12935 20156
rect 12935 20100 12939 20156
rect 12875 20096 12939 20100
rect 12955 20156 13019 20160
rect 12955 20100 12959 20156
rect 12959 20100 13015 20156
rect 13015 20100 13019 20156
rect 12955 20096 13019 20100
rect 20557 20156 20621 20160
rect 20557 20100 20561 20156
rect 20561 20100 20617 20156
rect 20617 20100 20621 20156
rect 20557 20096 20621 20100
rect 20637 20156 20701 20160
rect 20637 20100 20641 20156
rect 20641 20100 20697 20156
rect 20697 20100 20701 20156
rect 20637 20096 20701 20100
rect 20717 20156 20781 20160
rect 20717 20100 20721 20156
rect 20721 20100 20777 20156
rect 20777 20100 20781 20156
rect 20717 20096 20781 20100
rect 20797 20156 20861 20160
rect 20797 20100 20801 20156
rect 20801 20100 20857 20156
rect 20857 20100 20861 20156
rect 20797 20096 20861 20100
rect 28399 20156 28463 20160
rect 28399 20100 28403 20156
rect 28403 20100 28459 20156
rect 28459 20100 28463 20156
rect 28399 20096 28463 20100
rect 28479 20156 28543 20160
rect 28479 20100 28483 20156
rect 28483 20100 28539 20156
rect 28539 20100 28543 20156
rect 28479 20096 28543 20100
rect 28559 20156 28623 20160
rect 28559 20100 28563 20156
rect 28563 20100 28619 20156
rect 28619 20100 28623 20156
rect 28559 20096 28623 20100
rect 28639 20156 28703 20160
rect 28639 20100 28643 20156
rect 28643 20100 28699 20156
rect 28699 20100 28703 20156
rect 28639 20096 28703 20100
rect 8794 19612 8858 19616
rect 8794 19556 8798 19612
rect 8798 19556 8854 19612
rect 8854 19556 8858 19612
rect 8794 19552 8858 19556
rect 8874 19612 8938 19616
rect 8874 19556 8878 19612
rect 8878 19556 8934 19612
rect 8934 19556 8938 19612
rect 8874 19552 8938 19556
rect 8954 19612 9018 19616
rect 8954 19556 8958 19612
rect 8958 19556 9014 19612
rect 9014 19556 9018 19612
rect 8954 19552 9018 19556
rect 9034 19612 9098 19616
rect 9034 19556 9038 19612
rect 9038 19556 9094 19612
rect 9094 19556 9098 19612
rect 9034 19552 9098 19556
rect 16636 19612 16700 19616
rect 16636 19556 16640 19612
rect 16640 19556 16696 19612
rect 16696 19556 16700 19612
rect 16636 19552 16700 19556
rect 16716 19612 16780 19616
rect 16716 19556 16720 19612
rect 16720 19556 16776 19612
rect 16776 19556 16780 19612
rect 16716 19552 16780 19556
rect 16796 19612 16860 19616
rect 16796 19556 16800 19612
rect 16800 19556 16856 19612
rect 16856 19556 16860 19612
rect 16796 19552 16860 19556
rect 16876 19612 16940 19616
rect 16876 19556 16880 19612
rect 16880 19556 16936 19612
rect 16936 19556 16940 19612
rect 16876 19552 16940 19556
rect 24478 19612 24542 19616
rect 24478 19556 24482 19612
rect 24482 19556 24538 19612
rect 24538 19556 24542 19612
rect 24478 19552 24542 19556
rect 24558 19612 24622 19616
rect 24558 19556 24562 19612
rect 24562 19556 24618 19612
rect 24618 19556 24622 19612
rect 24558 19552 24622 19556
rect 24638 19612 24702 19616
rect 24638 19556 24642 19612
rect 24642 19556 24698 19612
rect 24698 19556 24702 19612
rect 24638 19552 24702 19556
rect 24718 19612 24782 19616
rect 24718 19556 24722 19612
rect 24722 19556 24778 19612
rect 24778 19556 24782 19612
rect 24718 19552 24782 19556
rect 32320 19612 32384 19616
rect 32320 19556 32324 19612
rect 32324 19556 32380 19612
rect 32380 19556 32384 19612
rect 32320 19552 32384 19556
rect 32400 19612 32464 19616
rect 32400 19556 32404 19612
rect 32404 19556 32460 19612
rect 32460 19556 32464 19612
rect 32400 19552 32464 19556
rect 32480 19612 32544 19616
rect 32480 19556 32484 19612
rect 32484 19556 32540 19612
rect 32540 19556 32544 19612
rect 32480 19552 32544 19556
rect 32560 19612 32624 19616
rect 32560 19556 32564 19612
rect 32564 19556 32620 19612
rect 32620 19556 32624 19612
rect 32560 19552 32624 19556
rect 2268 19484 2332 19548
rect 18460 19484 18524 19548
rect 13676 19408 13740 19412
rect 13676 19352 13726 19408
rect 13726 19352 13740 19408
rect 13676 19348 13740 19352
rect 4873 19068 4937 19072
rect 4873 19012 4877 19068
rect 4877 19012 4933 19068
rect 4933 19012 4937 19068
rect 4873 19008 4937 19012
rect 4953 19068 5017 19072
rect 4953 19012 4957 19068
rect 4957 19012 5013 19068
rect 5013 19012 5017 19068
rect 4953 19008 5017 19012
rect 5033 19068 5097 19072
rect 5033 19012 5037 19068
rect 5037 19012 5093 19068
rect 5093 19012 5097 19068
rect 5033 19008 5097 19012
rect 5113 19068 5177 19072
rect 5113 19012 5117 19068
rect 5117 19012 5173 19068
rect 5173 19012 5177 19068
rect 5113 19008 5177 19012
rect 12715 19068 12779 19072
rect 12715 19012 12719 19068
rect 12719 19012 12775 19068
rect 12775 19012 12779 19068
rect 12715 19008 12779 19012
rect 12795 19068 12859 19072
rect 12795 19012 12799 19068
rect 12799 19012 12855 19068
rect 12855 19012 12859 19068
rect 12795 19008 12859 19012
rect 12875 19068 12939 19072
rect 12875 19012 12879 19068
rect 12879 19012 12935 19068
rect 12935 19012 12939 19068
rect 12875 19008 12939 19012
rect 12955 19068 13019 19072
rect 12955 19012 12959 19068
rect 12959 19012 13015 19068
rect 13015 19012 13019 19068
rect 12955 19008 13019 19012
rect 20557 19068 20621 19072
rect 20557 19012 20561 19068
rect 20561 19012 20617 19068
rect 20617 19012 20621 19068
rect 20557 19008 20621 19012
rect 20637 19068 20701 19072
rect 20637 19012 20641 19068
rect 20641 19012 20697 19068
rect 20697 19012 20701 19068
rect 20637 19008 20701 19012
rect 20717 19068 20781 19072
rect 20717 19012 20721 19068
rect 20721 19012 20777 19068
rect 20777 19012 20781 19068
rect 20717 19008 20781 19012
rect 20797 19068 20861 19072
rect 20797 19012 20801 19068
rect 20801 19012 20857 19068
rect 20857 19012 20861 19068
rect 20797 19008 20861 19012
rect 28399 19068 28463 19072
rect 28399 19012 28403 19068
rect 28403 19012 28459 19068
rect 28459 19012 28463 19068
rect 28399 19008 28463 19012
rect 28479 19068 28543 19072
rect 28479 19012 28483 19068
rect 28483 19012 28539 19068
rect 28539 19012 28543 19068
rect 28479 19008 28543 19012
rect 28559 19068 28623 19072
rect 28559 19012 28563 19068
rect 28563 19012 28619 19068
rect 28619 19012 28623 19068
rect 28559 19008 28623 19012
rect 28639 19068 28703 19072
rect 28639 19012 28643 19068
rect 28643 19012 28699 19068
rect 28699 19012 28703 19068
rect 28639 19008 28703 19012
rect 8794 18524 8858 18528
rect 8794 18468 8798 18524
rect 8798 18468 8854 18524
rect 8854 18468 8858 18524
rect 8794 18464 8858 18468
rect 8874 18524 8938 18528
rect 8874 18468 8878 18524
rect 8878 18468 8934 18524
rect 8934 18468 8938 18524
rect 8874 18464 8938 18468
rect 8954 18524 9018 18528
rect 8954 18468 8958 18524
rect 8958 18468 9014 18524
rect 9014 18468 9018 18524
rect 8954 18464 9018 18468
rect 9034 18524 9098 18528
rect 9034 18468 9038 18524
rect 9038 18468 9094 18524
rect 9094 18468 9098 18524
rect 9034 18464 9098 18468
rect 16636 18524 16700 18528
rect 16636 18468 16640 18524
rect 16640 18468 16696 18524
rect 16696 18468 16700 18524
rect 16636 18464 16700 18468
rect 16716 18524 16780 18528
rect 16716 18468 16720 18524
rect 16720 18468 16776 18524
rect 16776 18468 16780 18524
rect 16716 18464 16780 18468
rect 16796 18524 16860 18528
rect 16796 18468 16800 18524
rect 16800 18468 16856 18524
rect 16856 18468 16860 18524
rect 16796 18464 16860 18468
rect 16876 18524 16940 18528
rect 16876 18468 16880 18524
rect 16880 18468 16936 18524
rect 16936 18468 16940 18524
rect 16876 18464 16940 18468
rect 24478 18524 24542 18528
rect 24478 18468 24482 18524
rect 24482 18468 24538 18524
rect 24538 18468 24542 18524
rect 24478 18464 24542 18468
rect 24558 18524 24622 18528
rect 24558 18468 24562 18524
rect 24562 18468 24618 18524
rect 24618 18468 24622 18524
rect 24558 18464 24622 18468
rect 24638 18524 24702 18528
rect 24638 18468 24642 18524
rect 24642 18468 24698 18524
rect 24698 18468 24702 18524
rect 24638 18464 24702 18468
rect 24718 18524 24782 18528
rect 24718 18468 24722 18524
rect 24722 18468 24778 18524
rect 24778 18468 24782 18524
rect 24718 18464 24782 18468
rect 32320 18524 32384 18528
rect 32320 18468 32324 18524
rect 32324 18468 32380 18524
rect 32380 18468 32384 18524
rect 32320 18464 32384 18468
rect 32400 18524 32464 18528
rect 32400 18468 32404 18524
rect 32404 18468 32460 18524
rect 32460 18468 32464 18524
rect 32400 18464 32464 18468
rect 32480 18524 32544 18528
rect 32480 18468 32484 18524
rect 32484 18468 32540 18524
rect 32540 18468 32544 18524
rect 32480 18464 32544 18468
rect 32560 18524 32624 18528
rect 32560 18468 32564 18524
rect 32564 18468 32620 18524
rect 32620 18468 32624 18524
rect 32560 18464 32624 18468
rect 4873 17980 4937 17984
rect 4873 17924 4877 17980
rect 4877 17924 4933 17980
rect 4933 17924 4937 17980
rect 4873 17920 4937 17924
rect 4953 17980 5017 17984
rect 4953 17924 4957 17980
rect 4957 17924 5013 17980
rect 5013 17924 5017 17980
rect 4953 17920 5017 17924
rect 5033 17980 5097 17984
rect 5033 17924 5037 17980
rect 5037 17924 5093 17980
rect 5093 17924 5097 17980
rect 5033 17920 5097 17924
rect 5113 17980 5177 17984
rect 5113 17924 5117 17980
rect 5117 17924 5173 17980
rect 5173 17924 5177 17980
rect 5113 17920 5177 17924
rect 12715 17980 12779 17984
rect 12715 17924 12719 17980
rect 12719 17924 12775 17980
rect 12775 17924 12779 17980
rect 12715 17920 12779 17924
rect 12795 17980 12859 17984
rect 12795 17924 12799 17980
rect 12799 17924 12855 17980
rect 12855 17924 12859 17980
rect 12795 17920 12859 17924
rect 12875 17980 12939 17984
rect 12875 17924 12879 17980
rect 12879 17924 12935 17980
rect 12935 17924 12939 17980
rect 12875 17920 12939 17924
rect 12955 17980 13019 17984
rect 12955 17924 12959 17980
rect 12959 17924 13015 17980
rect 13015 17924 13019 17980
rect 12955 17920 13019 17924
rect 20557 17980 20621 17984
rect 20557 17924 20561 17980
rect 20561 17924 20617 17980
rect 20617 17924 20621 17980
rect 20557 17920 20621 17924
rect 20637 17980 20701 17984
rect 20637 17924 20641 17980
rect 20641 17924 20697 17980
rect 20697 17924 20701 17980
rect 20637 17920 20701 17924
rect 20717 17980 20781 17984
rect 20717 17924 20721 17980
rect 20721 17924 20777 17980
rect 20777 17924 20781 17980
rect 20717 17920 20781 17924
rect 20797 17980 20861 17984
rect 20797 17924 20801 17980
rect 20801 17924 20857 17980
rect 20857 17924 20861 17980
rect 20797 17920 20861 17924
rect 28399 17980 28463 17984
rect 28399 17924 28403 17980
rect 28403 17924 28459 17980
rect 28459 17924 28463 17980
rect 28399 17920 28463 17924
rect 28479 17980 28543 17984
rect 28479 17924 28483 17980
rect 28483 17924 28539 17980
rect 28539 17924 28543 17980
rect 28479 17920 28543 17924
rect 28559 17980 28623 17984
rect 28559 17924 28563 17980
rect 28563 17924 28619 17980
rect 28619 17924 28623 17980
rect 28559 17920 28623 17924
rect 28639 17980 28703 17984
rect 28639 17924 28643 17980
rect 28643 17924 28699 17980
rect 28699 17924 28703 17980
rect 28639 17920 28703 17924
rect 1532 17912 1596 17916
rect 1532 17856 1582 17912
rect 1582 17856 1596 17912
rect 1532 17852 1596 17856
rect 3740 17852 3804 17916
rect 31524 17852 31588 17916
rect 8794 17436 8858 17440
rect 8794 17380 8798 17436
rect 8798 17380 8854 17436
rect 8854 17380 8858 17436
rect 8794 17376 8858 17380
rect 8874 17436 8938 17440
rect 8874 17380 8878 17436
rect 8878 17380 8934 17436
rect 8934 17380 8938 17436
rect 8874 17376 8938 17380
rect 8954 17436 9018 17440
rect 8954 17380 8958 17436
rect 8958 17380 9014 17436
rect 9014 17380 9018 17436
rect 8954 17376 9018 17380
rect 9034 17436 9098 17440
rect 9034 17380 9038 17436
rect 9038 17380 9094 17436
rect 9094 17380 9098 17436
rect 9034 17376 9098 17380
rect 16636 17436 16700 17440
rect 16636 17380 16640 17436
rect 16640 17380 16696 17436
rect 16696 17380 16700 17436
rect 16636 17376 16700 17380
rect 16716 17436 16780 17440
rect 16716 17380 16720 17436
rect 16720 17380 16776 17436
rect 16776 17380 16780 17436
rect 16716 17376 16780 17380
rect 16796 17436 16860 17440
rect 16796 17380 16800 17436
rect 16800 17380 16856 17436
rect 16856 17380 16860 17436
rect 16796 17376 16860 17380
rect 16876 17436 16940 17440
rect 16876 17380 16880 17436
rect 16880 17380 16936 17436
rect 16936 17380 16940 17436
rect 16876 17376 16940 17380
rect 24478 17436 24542 17440
rect 24478 17380 24482 17436
rect 24482 17380 24538 17436
rect 24538 17380 24542 17436
rect 24478 17376 24542 17380
rect 24558 17436 24622 17440
rect 24558 17380 24562 17436
rect 24562 17380 24618 17436
rect 24618 17380 24622 17436
rect 24558 17376 24622 17380
rect 24638 17436 24702 17440
rect 24638 17380 24642 17436
rect 24642 17380 24698 17436
rect 24698 17380 24702 17436
rect 24638 17376 24702 17380
rect 24718 17436 24782 17440
rect 24718 17380 24722 17436
rect 24722 17380 24778 17436
rect 24778 17380 24782 17436
rect 24718 17376 24782 17380
rect 32320 17436 32384 17440
rect 32320 17380 32324 17436
rect 32324 17380 32380 17436
rect 32380 17380 32384 17436
rect 32320 17376 32384 17380
rect 32400 17436 32464 17440
rect 32400 17380 32404 17436
rect 32404 17380 32460 17436
rect 32460 17380 32464 17436
rect 32400 17376 32464 17380
rect 32480 17436 32544 17440
rect 32480 17380 32484 17436
rect 32484 17380 32540 17436
rect 32540 17380 32544 17436
rect 32480 17376 32544 17380
rect 32560 17436 32624 17440
rect 32560 17380 32564 17436
rect 32564 17380 32620 17436
rect 32620 17380 32624 17436
rect 32560 17376 32624 17380
rect 30236 16960 30300 16964
rect 30236 16904 30286 16960
rect 30286 16904 30300 16960
rect 30236 16900 30300 16904
rect 4873 16892 4937 16896
rect 4873 16836 4877 16892
rect 4877 16836 4933 16892
rect 4933 16836 4937 16892
rect 4873 16832 4937 16836
rect 4953 16892 5017 16896
rect 4953 16836 4957 16892
rect 4957 16836 5013 16892
rect 5013 16836 5017 16892
rect 4953 16832 5017 16836
rect 5033 16892 5097 16896
rect 5033 16836 5037 16892
rect 5037 16836 5093 16892
rect 5093 16836 5097 16892
rect 5033 16832 5097 16836
rect 5113 16892 5177 16896
rect 5113 16836 5117 16892
rect 5117 16836 5173 16892
rect 5173 16836 5177 16892
rect 5113 16832 5177 16836
rect 12715 16892 12779 16896
rect 12715 16836 12719 16892
rect 12719 16836 12775 16892
rect 12775 16836 12779 16892
rect 12715 16832 12779 16836
rect 12795 16892 12859 16896
rect 12795 16836 12799 16892
rect 12799 16836 12855 16892
rect 12855 16836 12859 16892
rect 12795 16832 12859 16836
rect 12875 16892 12939 16896
rect 12875 16836 12879 16892
rect 12879 16836 12935 16892
rect 12935 16836 12939 16892
rect 12875 16832 12939 16836
rect 12955 16892 13019 16896
rect 12955 16836 12959 16892
rect 12959 16836 13015 16892
rect 13015 16836 13019 16892
rect 12955 16832 13019 16836
rect 20557 16892 20621 16896
rect 20557 16836 20561 16892
rect 20561 16836 20617 16892
rect 20617 16836 20621 16892
rect 20557 16832 20621 16836
rect 20637 16892 20701 16896
rect 20637 16836 20641 16892
rect 20641 16836 20697 16892
rect 20697 16836 20701 16892
rect 20637 16832 20701 16836
rect 20717 16892 20781 16896
rect 20717 16836 20721 16892
rect 20721 16836 20777 16892
rect 20777 16836 20781 16892
rect 20717 16832 20781 16836
rect 20797 16892 20861 16896
rect 20797 16836 20801 16892
rect 20801 16836 20857 16892
rect 20857 16836 20861 16892
rect 20797 16832 20861 16836
rect 28399 16892 28463 16896
rect 28399 16836 28403 16892
rect 28403 16836 28459 16892
rect 28459 16836 28463 16892
rect 28399 16832 28463 16836
rect 28479 16892 28543 16896
rect 28479 16836 28483 16892
rect 28483 16836 28539 16892
rect 28539 16836 28543 16892
rect 28479 16832 28543 16836
rect 28559 16892 28623 16896
rect 28559 16836 28563 16892
rect 28563 16836 28619 16892
rect 28619 16836 28623 16892
rect 28559 16832 28623 16836
rect 28639 16892 28703 16896
rect 28639 16836 28643 16892
rect 28643 16836 28699 16892
rect 28699 16836 28703 16892
rect 28639 16832 28703 16836
rect 8794 16348 8858 16352
rect 8794 16292 8798 16348
rect 8798 16292 8854 16348
rect 8854 16292 8858 16348
rect 8794 16288 8858 16292
rect 8874 16348 8938 16352
rect 8874 16292 8878 16348
rect 8878 16292 8934 16348
rect 8934 16292 8938 16348
rect 8874 16288 8938 16292
rect 8954 16348 9018 16352
rect 8954 16292 8958 16348
rect 8958 16292 9014 16348
rect 9014 16292 9018 16348
rect 8954 16288 9018 16292
rect 9034 16348 9098 16352
rect 9034 16292 9038 16348
rect 9038 16292 9094 16348
rect 9094 16292 9098 16348
rect 9034 16288 9098 16292
rect 16636 16348 16700 16352
rect 16636 16292 16640 16348
rect 16640 16292 16696 16348
rect 16696 16292 16700 16348
rect 16636 16288 16700 16292
rect 16716 16348 16780 16352
rect 16716 16292 16720 16348
rect 16720 16292 16776 16348
rect 16776 16292 16780 16348
rect 16716 16288 16780 16292
rect 16796 16348 16860 16352
rect 16796 16292 16800 16348
rect 16800 16292 16856 16348
rect 16856 16292 16860 16348
rect 16796 16288 16860 16292
rect 16876 16348 16940 16352
rect 16876 16292 16880 16348
rect 16880 16292 16936 16348
rect 16936 16292 16940 16348
rect 16876 16288 16940 16292
rect 24478 16348 24542 16352
rect 24478 16292 24482 16348
rect 24482 16292 24538 16348
rect 24538 16292 24542 16348
rect 24478 16288 24542 16292
rect 24558 16348 24622 16352
rect 24558 16292 24562 16348
rect 24562 16292 24618 16348
rect 24618 16292 24622 16348
rect 24558 16288 24622 16292
rect 24638 16348 24702 16352
rect 24638 16292 24642 16348
rect 24642 16292 24698 16348
rect 24698 16292 24702 16348
rect 24638 16288 24702 16292
rect 24718 16348 24782 16352
rect 24718 16292 24722 16348
rect 24722 16292 24778 16348
rect 24778 16292 24782 16348
rect 24718 16288 24782 16292
rect 32320 16348 32384 16352
rect 32320 16292 32324 16348
rect 32324 16292 32380 16348
rect 32380 16292 32384 16348
rect 32320 16288 32384 16292
rect 32400 16348 32464 16352
rect 32400 16292 32404 16348
rect 32404 16292 32460 16348
rect 32460 16292 32464 16348
rect 32400 16288 32464 16292
rect 32480 16348 32544 16352
rect 32480 16292 32484 16348
rect 32484 16292 32540 16348
rect 32540 16292 32544 16348
rect 32480 16288 32544 16292
rect 32560 16348 32624 16352
rect 32560 16292 32564 16348
rect 32564 16292 32620 16348
rect 32620 16292 32624 16348
rect 32560 16288 32624 16292
rect 4873 15804 4937 15808
rect 4873 15748 4877 15804
rect 4877 15748 4933 15804
rect 4933 15748 4937 15804
rect 4873 15744 4937 15748
rect 4953 15804 5017 15808
rect 4953 15748 4957 15804
rect 4957 15748 5013 15804
rect 5013 15748 5017 15804
rect 4953 15744 5017 15748
rect 5033 15804 5097 15808
rect 5033 15748 5037 15804
rect 5037 15748 5093 15804
rect 5093 15748 5097 15804
rect 5033 15744 5097 15748
rect 5113 15804 5177 15808
rect 5113 15748 5117 15804
rect 5117 15748 5173 15804
rect 5173 15748 5177 15804
rect 5113 15744 5177 15748
rect 12715 15804 12779 15808
rect 12715 15748 12719 15804
rect 12719 15748 12775 15804
rect 12775 15748 12779 15804
rect 12715 15744 12779 15748
rect 12795 15804 12859 15808
rect 12795 15748 12799 15804
rect 12799 15748 12855 15804
rect 12855 15748 12859 15804
rect 12795 15744 12859 15748
rect 12875 15804 12939 15808
rect 12875 15748 12879 15804
rect 12879 15748 12935 15804
rect 12935 15748 12939 15804
rect 12875 15744 12939 15748
rect 12955 15804 13019 15808
rect 12955 15748 12959 15804
rect 12959 15748 13015 15804
rect 13015 15748 13019 15804
rect 12955 15744 13019 15748
rect 20557 15804 20621 15808
rect 20557 15748 20561 15804
rect 20561 15748 20617 15804
rect 20617 15748 20621 15804
rect 20557 15744 20621 15748
rect 20637 15804 20701 15808
rect 20637 15748 20641 15804
rect 20641 15748 20697 15804
rect 20697 15748 20701 15804
rect 20637 15744 20701 15748
rect 20717 15804 20781 15808
rect 20717 15748 20721 15804
rect 20721 15748 20777 15804
rect 20777 15748 20781 15804
rect 20717 15744 20781 15748
rect 20797 15804 20861 15808
rect 20797 15748 20801 15804
rect 20801 15748 20857 15804
rect 20857 15748 20861 15804
rect 20797 15744 20861 15748
rect 28399 15804 28463 15808
rect 28399 15748 28403 15804
rect 28403 15748 28459 15804
rect 28459 15748 28463 15804
rect 28399 15744 28463 15748
rect 28479 15804 28543 15808
rect 28479 15748 28483 15804
rect 28483 15748 28539 15804
rect 28539 15748 28543 15804
rect 28479 15744 28543 15748
rect 28559 15804 28623 15808
rect 28559 15748 28563 15804
rect 28563 15748 28619 15804
rect 28619 15748 28623 15804
rect 28559 15744 28623 15748
rect 28639 15804 28703 15808
rect 28639 15748 28643 15804
rect 28643 15748 28699 15804
rect 28699 15748 28703 15804
rect 28639 15744 28703 15748
rect 8794 15260 8858 15264
rect 8794 15204 8798 15260
rect 8798 15204 8854 15260
rect 8854 15204 8858 15260
rect 8794 15200 8858 15204
rect 8874 15260 8938 15264
rect 8874 15204 8878 15260
rect 8878 15204 8934 15260
rect 8934 15204 8938 15260
rect 8874 15200 8938 15204
rect 8954 15260 9018 15264
rect 8954 15204 8958 15260
rect 8958 15204 9014 15260
rect 9014 15204 9018 15260
rect 8954 15200 9018 15204
rect 9034 15260 9098 15264
rect 9034 15204 9038 15260
rect 9038 15204 9094 15260
rect 9094 15204 9098 15260
rect 9034 15200 9098 15204
rect 16636 15260 16700 15264
rect 16636 15204 16640 15260
rect 16640 15204 16696 15260
rect 16696 15204 16700 15260
rect 16636 15200 16700 15204
rect 16716 15260 16780 15264
rect 16716 15204 16720 15260
rect 16720 15204 16776 15260
rect 16776 15204 16780 15260
rect 16716 15200 16780 15204
rect 16796 15260 16860 15264
rect 16796 15204 16800 15260
rect 16800 15204 16856 15260
rect 16856 15204 16860 15260
rect 16796 15200 16860 15204
rect 16876 15260 16940 15264
rect 16876 15204 16880 15260
rect 16880 15204 16936 15260
rect 16936 15204 16940 15260
rect 16876 15200 16940 15204
rect 24478 15260 24542 15264
rect 24478 15204 24482 15260
rect 24482 15204 24538 15260
rect 24538 15204 24542 15260
rect 24478 15200 24542 15204
rect 24558 15260 24622 15264
rect 24558 15204 24562 15260
rect 24562 15204 24618 15260
rect 24618 15204 24622 15260
rect 24558 15200 24622 15204
rect 24638 15260 24702 15264
rect 24638 15204 24642 15260
rect 24642 15204 24698 15260
rect 24698 15204 24702 15260
rect 24638 15200 24702 15204
rect 24718 15260 24782 15264
rect 24718 15204 24722 15260
rect 24722 15204 24778 15260
rect 24778 15204 24782 15260
rect 24718 15200 24782 15204
rect 32320 15260 32384 15264
rect 32320 15204 32324 15260
rect 32324 15204 32380 15260
rect 32380 15204 32384 15260
rect 32320 15200 32384 15204
rect 32400 15260 32464 15264
rect 32400 15204 32404 15260
rect 32404 15204 32460 15260
rect 32460 15204 32464 15260
rect 32400 15200 32464 15204
rect 32480 15260 32544 15264
rect 32480 15204 32484 15260
rect 32484 15204 32540 15260
rect 32540 15204 32544 15260
rect 32480 15200 32544 15204
rect 32560 15260 32624 15264
rect 32560 15204 32564 15260
rect 32564 15204 32620 15260
rect 32620 15204 32624 15260
rect 32560 15200 32624 15204
rect 4873 14716 4937 14720
rect 4873 14660 4877 14716
rect 4877 14660 4933 14716
rect 4933 14660 4937 14716
rect 4873 14656 4937 14660
rect 4953 14716 5017 14720
rect 4953 14660 4957 14716
rect 4957 14660 5013 14716
rect 5013 14660 5017 14716
rect 4953 14656 5017 14660
rect 5033 14716 5097 14720
rect 5033 14660 5037 14716
rect 5037 14660 5093 14716
rect 5093 14660 5097 14716
rect 5033 14656 5097 14660
rect 5113 14716 5177 14720
rect 5113 14660 5117 14716
rect 5117 14660 5173 14716
rect 5173 14660 5177 14716
rect 5113 14656 5177 14660
rect 12715 14716 12779 14720
rect 12715 14660 12719 14716
rect 12719 14660 12775 14716
rect 12775 14660 12779 14716
rect 12715 14656 12779 14660
rect 12795 14716 12859 14720
rect 12795 14660 12799 14716
rect 12799 14660 12855 14716
rect 12855 14660 12859 14716
rect 12795 14656 12859 14660
rect 12875 14716 12939 14720
rect 12875 14660 12879 14716
rect 12879 14660 12935 14716
rect 12935 14660 12939 14716
rect 12875 14656 12939 14660
rect 12955 14716 13019 14720
rect 12955 14660 12959 14716
rect 12959 14660 13015 14716
rect 13015 14660 13019 14716
rect 12955 14656 13019 14660
rect 20557 14716 20621 14720
rect 20557 14660 20561 14716
rect 20561 14660 20617 14716
rect 20617 14660 20621 14716
rect 20557 14656 20621 14660
rect 20637 14716 20701 14720
rect 20637 14660 20641 14716
rect 20641 14660 20697 14716
rect 20697 14660 20701 14716
rect 20637 14656 20701 14660
rect 20717 14716 20781 14720
rect 20717 14660 20721 14716
rect 20721 14660 20777 14716
rect 20777 14660 20781 14716
rect 20717 14656 20781 14660
rect 20797 14716 20861 14720
rect 20797 14660 20801 14716
rect 20801 14660 20857 14716
rect 20857 14660 20861 14716
rect 20797 14656 20861 14660
rect 28399 14716 28463 14720
rect 28399 14660 28403 14716
rect 28403 14660 28459 14716
rect 28459 14660 28463 14716
rect 28399 14656 28463 14660
rect 28479 14716 28543 14720
rect 28479 14660 28483 14716
rect 28483 14660 28539 14716
rect 28539 14660 28543 14716
rect 28479 14656 28543 14660
rect 28559 14716 28623 14720
rect 28559 14660 28563 14716
rect 28563 14660 28619 14716
rect 28619 14660 28623 14716
rect 28559 14656 28623 14660
rect 28639 14716 28703 14720
rect 28639 14660 28643 14716
rect 28643 14660 28699 14716
rect 28699 14660 28703 14716
rect 28639 14656 28703 14660
rect 8794 14172 8858 14176
rect 8794 14116 8798 14172
rect 8798 14116 8854 14172
rect 8854 14116 8858 14172
rect 8794 14112 8858 14116
rect 8874 14172 8938 14176
rect 8874 14116 8878 14172
rect 8878 14116 8934 14172
rect 8934 14116 8938 14172
rect 8874 14112 8938 14116
rect 8954 14172 9018 14176
rect 8954 14116 8958 14172
rect 8958 14116 9014 14172
rect 9014 14116 9018 14172
rect 8954 14112 9018 14116
rect 9034 14172 9098 14176
rect 9034 14116 9038 14172
rect 9038 14116 9094 14172
rect 9094 14116 9098 14172
rect 9034 14112 9098 14116
rect 16636 14172 16700 14176
rect 16636 14116 16640 14172
rect 16640 14116 16696 14172
rect 16696 14116 16700 14172
rect 16636 14112 16700 14116
rect 16716 14172 16780 14176
rect 16716 14116 16720 14172
rect 16720 14116 16776 14172
rect 16776 14116 16780 14172
rect 16716 14112 16780 14116
rect 16796 14172 16860 14176
rect 16796 14116 16800 14172
rect 16800 14116 16856 14172
rect 16856 14116 16860 14172
rect 16796 14112 16860 14116
rect 16876 14172 16940 14176
rect 16876 14116 16880 14172
rect 16880 14116 16936 14172
rect 16936 14116 16940 14172
rect 16876 14112 16940 14116
rect 24478 14172 24542 14176
rect 24478 14116 24482 14172
rect 24482 14116 24538 14172
rect 24538 14116 24542 14172
rect 24478 14112 24542 14116
rect 24558 14172 24622 14176
rect 24558 14116 24562 14172
rect 24562 14116 24618 14172
rect 24618 14116 24622 14172
rect 24558 14112 24622 14116
rect 24638 14172 24702 14176
rect 24638 14116 24642 14172
rect 24642 14116 24698 14172
rect 24698 14116 24702 14172
rect 24638 14112 24702 14116
rect 24718 14172 24782 14176
rect 24718 14116 24722 14172
rect 24722 14116 24778 14172
rect 24778 14116 24782 14172
rect 24718 14112 24782 14116
rect 32320 14172 32384 14176
rect 32320 14116 32324 14172
rect 32324 14116 32380 14172
rect 32380 14116 32384 14172
rect 32320 14112 32384 14116
rect 32400 14172 32464 14176
rect 32400 14116 32404 14172
rect 32404 14116 32460 14172
rect 32460 14116 32464 14172
rect 32400 14112 32464 14116
rect 32480 14172 32544 14176
rect 32480 14116 32484 14172
rect 32484 14116 32540 14172
rect 32540 14116 32544 14172
rect 32480 14112 32544 14116
rect 32560 14172 32624 14176
rect 32560 14116 32564 14172
rect 32564 14116 32620 14172
rect 32620 14116 32624 14172
rect 32560 14112 32624 14116
rect 4873 13628 4937 13632
rect 4873 13572 4877 13628
rect 4877 13572 4933 13628
rect 4933 13572 4937 13628
rect 4873 13568 4937 13572
rect 4953 13628 5017 13632
rect 4953 13572 4957 13628
rect 4957 13572 5013 13628
rect 5013 13572 5017 13628
rect 4953 13568 5017 13572
rect 5033 13628 5097 13632
rect 5033 13572 5037 13628
rect 5037 13572 5093 13628
rect 5093 13572 5097 13628
rect 5033 13568 5097 13572
rect 5113 13628 5177 13632
rect 5113 13572 5117 13628
rect 5117 13572 5173 13628
rect 5173 13572 5177 13628
rect 5113 13568 5177 13572
rect 12715 13628 12779 13632
rect 12715 13572 12719 13628
rect 12719 13572 12775 13628
rect 12775 13572 12779 13628
rect 12715 13568 12779 13572
rect 12795 13628 12859 13632
rect 12795 13572 12799 13628
rect 12799 13572 12855 13628
rect 12855 13572 12859 13628
rect 12795 13568 12859 13572
rect 12875 13628 12939 13632
rect 12875 13572 12879 13628
rect 12879 13572 12935 13628
rect 12935 13572 12939 13628
rect 12875 13568 12939 13572
rect 12955 13628 13019 13632
rect 12955 13572 12959 13628
rect 12959 13572 13015 13628
rect 13015 13572 13019 13628
rect 12955 13568 13019 13572
rect 20557 13628 20621 13632
rect 20557 13572 20561 13628
rect 20561 13572 20617 13628
rect 20617 13572 20621 13628
rect 20557 13568 20621 13572
rect 20637 13628 20701 13632
rect 20637 13572 20641 13628
rect 20641 13572 20697 13628
rect 20697 13572 20701 13628
rect 20637 13568 20701 13572
rect 20717 13628 20781 13632
rect 20717 13572 20721 13628
rect 20721 13572 20777 13628
rect 20777 13572 20781 13628
rect 20717 13568 20781 13572
rect 20797 13628 20861 13632
rect 20797 13572 20801 13628
rect 20801 13572 20857 13628
rect 20857 13572 20861 13628
rect 20797 13568 20861 13572
rect 28399 13628 28463 13632
rect 28399 13572 28403 13628
rect 28403 13572 28459 13628
rect 28459 13572 28463 13628
rect 28399 13568 28463 13572
rect 28479 13628 28543 13632
rect 28479 13572 28483 13628
rect 28483 13572 28539 13628
rect 28539 13572 28543 13628
rect 28479 13568 28543 13572
rect 28559 13628 28623 13632
rect 28559 13572 28563 13628
rect 28563 13572 28619 13628
rect 28619 13572 28623 13628
rect 28559 13568 28623 13572
rect 28639 13628 28703 13632
rect 28639 13572 28643 13628
rect 28643 13572 28699 13628
rect 28699 13572 28703 13628
rect 28639 13568 28703 13572
rect 8794 13084 8858 13088
rect 8794 13028 8798 13084
rect 8798 13028 8854 13084
rect 8854 13028 8858 13084
rect 8794 13024 8858 13028
rect 8874 13084 8938 13088
rect 8874 13028 8878 13084
rect 8878 13028 8934 13084
rect 8934 13028 8938 13084
rect 8874 13024 8938 13028
rect 8954 13084 9018 13088
rect 8954 13028 8958 13084
rect 8958 13028 9014 13084
rect 9014 13028 9018 13084
rect 8954 13024 9018 13028
rect 9034 13084 9098 13088
rect 9034 13028 9038 13084
rect 9038 13028 9094 13084
rect 9094 13028 9098 13084
rect 9034 13024 9098 13028
rect 16636 13084 16700 13088
rect 16636 13028 16640 13084
rect 16640 13028 16696 13084
rect 16696 13028 16700 13084
rect 16636 13024 16700 13028
rect 16716 13084 16780 13088
rect 16716 13028 16720 13084
rect 16720 13028 16776 13084
rect 16776 13028 16780 13084
rect 16716 13024 16780 13028
rect 16796 13084 16860 13088
rect 16796 13028 16800 13084
rect 16800 13028 16856 13084
rect 16856 13028 16860 13084
rect 16796 13024 16860 13028
rect 16876 13084 16940 13088
rect 16876 13028 16880 13084
rect 16880 13028 16936 13084
rect 16936 13028 16940 13084
rect 16876 13024 16940 13028
rect 24478 13084 24542 13088
rect 24478 13028 24482 13084
rect 24482 13028 24538 13084
rect 24538 13028 24542 13084
rect 24478 13024 24542 13028
rect 24558 13084 24622 13088
rect 24558 13028 24562 13084
rect 24562 13028 24618 13084
rect 24618 13028 24622 13084
rect 24558 13024 24622 13028
rect 24638 13084 24702 13088
rect 24638 13028 24642 13084
rect 24642 13028 24698 13084
rect 24698 13028 24702 13084
rect 24638 13024 24702 13028
rect 24718 13084 24782 13088
rect 24718 13028 24722 13084
rect 24722 13028 24778 13084
rect 24778 13028 24782 13084
rect 24718 13024 24782 13028
rect 32320 13084 32384 13088
rect 32320 13028 32324 13084
rect 32324 13028 32380 13084
rect 32380 13028 32384 13084
rect 32320 13024 32384 13028
rect 32400 13084 32464 13088
rect 32400 13028 32404 13084
rect 32404 13028 32460 13084
rect 32460 13028 32464 13084
rect 32400 13024 32464 13028
rect 32480 13084 32544 13088
rect 32480 13028 32484 13084
rect 32484 13028 32540 13084
rect 32540 13028 32544 13084
rect 32480 13024 32544 13028
rect 32560 13084 32624 13088
rect 32560 13028 32564 13084
rect 32564 13028 32620 13084
rect 32620 13028 32624 13084
rect 32560 13024 32624 13028
rect 4873 12540 4937 12544
rect 4873 12484 4877 12540
rect 4877 12484 4933 12540
rect 4933 12484 4937 12540
rect 4873 12480 4937 12484
rect 4953 12540 5017 12544
rect 4953 12484 4957 12540
rect 4957 12484 5013 12540
rect 5013 12484 5017 12540
rect 4953 12480 5017 12484
rect 5033 12540 5097 12544
rect 5033 12484 5037 12540
rect 5037 12484 5093 12540
rect 5093 12484 5097 12540
rect 5033 12480 5097 12484
rect 5113 12540 5177 12544
rect 5113 12484 5117 12540
rect 5117 12484 5173 12540
rect 5173 12484 5177 12540
rect 5113 12480 5177 12484
rect 12715 12540 12779 12544
rect 12715 12484 12719 12540
rect 12719 12484 12775 12540
rect 12775 12484 12779 12540
rect 12715 12480 12779 12484
rect 12795 12540 12859 12544
rect 12795 12484 12799 12540
rect 12799 12484 12855 12540
rect 12855 12484 12859 12540
rect 12795 12480 12859 12484
rect 12875 12540 12939 12544
rect 12875 12484 12879 12540
rect 12879 12484 12935 12540
rect 12935 12484 12939 12540
rect 12875 12480 12939 12484
rect 12955 12540 13019 12544
rect 12955 12484 12959 12540
rect 12959 12484 13015 12540
rect 13015 12484 13019 12540
rect 12955 12480 13019 12484
rect 20557 12540 20621 12544
rect 20557 12484 20561 12540
rect 20561 12484 20617 12540
rect 20617 12484 20621 12540
rect 20557 12480 20621 12484
rect 20637 12540 20701 12544
rect 20637 12484 20641 12540
rect 20641 12484 20697 12540
rect 20697 12484 20701 12540
rect 20637 12480 20701 12484
rect 20717 12540 20781 12544
rect 20717 12484 20721 12540
rect 20721 12484 20777 12540
rect 20777 12484 20781 12540
rect 20717 12480 20781 12484
rect 20797 12540 20861 12544
rect 20797 12484 20801 12540
rect 20801 12484 20857 12540
rect 20857 12484 20861 12540
rect 20797 12480 20861 12484
rect 28399 12540 28463 12544
rect 28399 12484 28403 12540
rect 28403 12484 28459 12540
rect 28459 12484 28463 12540
rect 28399 12480 28463 12484
rect 28479 12540 28543 12544
rect 28479 12484 28483 12540
rect 28483 12484 28539 12540
rect 28539 12484 28543 12540
rect 28479 12480 28543 12484
rect 28559 12540 28623 12544
rect 28559 12484 28563 12540
rect 28563 12484 28619 12540
rect 28619 12484 28623 12540
rect 28559 12480 28623 12484
rect 28639 12540 28703 12544
rect 28639 12484 28643 12540
rect 28643 12484 28699 12540
rect 28699 12484 28703 12540
rect 28639 12480 28703 12484
rect 13676 12276 13740 12340
rect 8794 11996 8858 12000
rect 8794 11940 8798 11996
rect 8798 11940 8854 11996
rect 8854 11940 8858 11996
rect 8794 11936 8858 11940
rect 8874 11996 8938 12000
rect 8874 11940 8878 11996
rect 8878 11940 8934 11996
rect 8934 11940 8938 11996
rect 8874 11936 8938 11940
rect 8954 11996 9018 12000
rect 8954 11940 8958 11996
rect 8958 11940 9014 11996
rect 9014 11940 9018 11996
rect 8954 11936 9018 11940
rect 9034 11996 9098 12000
rect 9034 11940 9038 11996
rect 9038 11940 9094 11996
rect 9094 11940 9098 11996
rect 9034 11936 9098 11940
rect 16636 11996 16700 12000
rect 16636 11940 16640 11996
rect 16640 11940 16696 11996
rect 16696 11940 16700 11996
rect 16636 11936 16700 11940
rect 16716 11996 16780 12000
rect 16716 11940 16720 11996
rect 16720 11940 16776 11996
rect 16776 11940 16780 11996
rect 16716 11936 16780 11940
rect 16796 11996 16860 12000
rect 16796 11940 16800 11996
rect 16800 11940 16856 11996
rect 16856 11940 16860 11996
rect 16796 11936 16860 11940
rect 16876 11996 16940 12000
rect 16876 11940 16880 11996
rect 16880 11940 16936 11996
rect 16936 11940 16940 11996
rect 16876 11936 16940 11940
rect 24478 11996 24542 12000
rect 24478 11940 24482 11996
rect 24482 11940 24538 11996
rect 24538 11940 24542 11996
rect 24478 11936 24542 11940
rect 24558 11996 24622 12000
rect 24558 11940 24562 11996
rect 24562 11940 24618 11996
rect 24618 11940 24622 11996
rect 24558 11936 24622 11940
rect 24638 11996 24702 12000
rect 24638 11940 24642 11996
rect 24642 11940 24698 11996
rect 24698 11940 24702 11996
rect 24638 11936 24702 11940
rect 24718 11996 24782 12000
rect 24718 11940 24722 11996
rect 24722 11940 24778 11996
rect 24778 11940 24782 11996
rect 24718 11936 24782 11940
rect 32320 11996 32384 12000
rect 32320 11940 32324 11996
rect 32324 11940 32380 11996
rect 32380 11940 32384 11996
rect 32320 11936 32384 11940
rect 32400 11996 32464 12000
rect 32400 11940 32404 11996
rect 32404 11940 32460 11996
rect 32460 11940 32464 11996
rect 32400 11936 32464 11940
rect 32480 11996 32544 12000
rect 32480 11940 32484 11996
rect 32484 11940 32540 11996
rect 32540 11940 32544 11996
rect 32480 11936 32544 11940
rect 32560 11996 32624 12000
rect 32560 11940 32564 11996
rect 32564 11940 32620 11996
rect 32620 11940 32624 11996
rect 32560 11936 32624 11940
rect 4873 11452 4937 11456
rect 4873 11396 4877 11452
rect 4877 11396 4933 11452
rect 4933 11396 4937 11452
rect 4873 11392 4937 11396
rect 4953 11452 5017 11456
rect 4953 11396 4957 11452
rect 4957 11396 5013 11452
rect 5013 11396 5017 11452
rect 4953 11392 5017 11396
rect 5033 11452 5097 11456
rect 5033 11396 5037 11452
rect 5037 11396 5093 11452
rect 5093 11396 5097 11452
rect 5033 11392 5097 11396
rect 5113 11452 5177 11456
rect 5113 11396 5117 11452
rect 5117 11396 5173 11452
rect 5173 11396 5177 11452
rect 5113 11392 5177 11396
rect 12715 11452 12779 11456
rect 12715 11396 12719 11452
rect 12719 11396 12775 11452
rect 12775 11396 12779 11452
rect 12715 11392 12779 11396
rect 12795 11452 12859 11456
rect 12795 11396 12799 11452
rect 12799 11396 12855 11452
rect 12855 11396 12859 11452
rect 12795 11392 12859 11396
rect 12875 11452 12939 11456
rect 12875 11396 12879 11452
rect 12879 11396 12935 11452
rect 12935 11396 12939 11452
rect 12875 11392 12939 11396
rect 12955 11452 13019 11456
rect 12955 11396 12959 11452
rect 12959 11396 13015 11452
rect 13015 11396 13019 11452
rect 12955 11392 13019 11396
rect 20557 11452 20621 11456
rect 20557 11396 20561 11452
rect 20561 11396 20617 11452
rect 20617 11396 20621 11452
rect 20557 11392 20621 11396
rect 20637 11452 20701 11456
rect 20637 11396 20641 11452
rect 20641 11396 20697 11452
rect 20697 11396 20701 11452
rect 20637 11392 20701 11396
rect 20717 11452 20781 11456
rect 20717 11396 20721 11452
rect 20721 11396 20777 11452
rect 20777 11396 20781 11452
rect 20717 11392 20781 11396
rect 20797 11452 20861 11456
rect 20797 11396 20801 11452
rect 20801 11396 20857 11452
rect 20857 11396 20861 11452
rect 20797 11392 20861 11396
rect 28399 11452 28463 11456
rect 28399 11396 28403 11452
rect 28403 11396 28459 11452
rect 28459 11396 28463 11452
rect 28399 11392 28463 11396
rect 28479 11452 28543 11456
rect 28479 11396 28483 11452
rect 28483 11396 28539 11452
rect 28539 11396 28543 11452
rect 28479 11392 28543 11396
rect 28559 11452 28623 11456
rect 28559 11396 28563 11452
rect 28563 11396 28619 11452
rect 28619 11396 28623 11452
rect 28559 11392 28623 11396
rect 28639 11452 28703 11456
rect 28639 11396 28643 11452
rect 28643 11396 28699 11452
rect 28699 11396 28703 11452
rect 28639 11392 28703 11396
rect 8794 10908 8858 10912
rect 8794 10852 8798 10908
rect 8798 10852 8854 10908
rect 8854 10852 8858 10908
rect 8794 10848 8858 10852
rect 8874 10908 8938 10912
rect 8874 10852 8878 10908
rect 8878 10852 8934 10908
rect 8934 10852 8938 10908
rect 8874 10848 8938 10852
rect 8954 10908 9018 10912
rect 8954 10852 8958 10908
rect 8958 10852 9014 10908
rect 9014 10852 9018 10908
rect 8954 10848 9018 10852
rect 9034 10908 9098 10912
rect 9034 10852 9038 10908
rect 9038 10852 9094 10908
rect 9094 10852 9098 10908
rect 9034 10848 9098 10852
rect 16636 10908 16700 10912
rect 16636 10852 16640 10908
rect 16640 10852 16696 10908
rect 16696 10852 16700 10908
rect 16636 10848 16700 10852
rect 16716 10908 16780 10912
rect 16716 10852 16720 10908
rect 16720 10852 16776 10908
rect 16776 10852 16780 10908
rect 16716 10848 16780 10852
rect 16796 10908 16860 10912
rect 16796 10852 16800 10908
rect 16800 10852 16856 10908
rect 16856 10852 16860 10908
rect 16796 10848 16860 10852
rect 16876 10908 16940 10912
rect 16876 10852 16880 10908
rect 16880 10852 16936 10908
rect 16936 10852 16940 10908
rect 16876 10848 16940 10852
rect 24478 10908 24542 10912
rect 24478 10852 24482 10908
rect 24482 10852 24538 10908
rect 24538 10852 24542 10908
rect 24478 10848 24542 10852
rect 24558 10908 24622 10912
rect 24558 10852 24562 10908
rect 24562 10852 24618 10908
rect 24618 10852 24622 10908
rect 24558 10848 24622 10852
rect 24638 10908 24702 10912
rect 24638 10852 24642 10908
rect 24642 10852 24698 10908
rect 24698 10852 24702 10908
rect 24638 10848 24702 10852
rect 24718 10908 24782 10912
rect 24718 10852 24722 10908
rect 24722 10852 24778 10908
rect 24778 10852 24782 10908
rect 24718 10848 24782 10852
rect 32320 10908 32384 10912
rect 32320 10852 32324 10908
rect 32324 10852 32380 10908
rect 32380 10852 32384 10908
rect 32320 10848 32384 10852
rect 32400 10908 32464 10912
rect 32400 10852 32404 10908
rect 32404 10852 32460 10908
rect 32460 10852 32464 10908
rect 32400 10848 32464 10852
rect 32480 10908 32544 10912
rect 32480 10852 32484 10908
rect 32484 10852 32540 10908
rect 32540 10852 32544 10908
rect 32480 10848 32544 10852
rect 32560 10908 32624 10912
rect 32560 10852 32564 10908
rect 32564 10852 32620 10908
rect 32620 10852 32624 10908
rect 32560 10848 32624 10852
rect 4873 10364 4937 10368
rect 4873 10308 4877 10364
rect 4877 10308 4933 10364
rect 4933 10308 4937 10364
rect 4873 10304 4937 10308
rect 4953 10364 5017 10368
rect 4953 10308 4957 10364
rect 4957 10308 5013 10364
rect 5013 10308 5017 10364
rect 4953 10304 5017 10308
rect 5033 10364 5097 10368
rect 5033 10308 5037 10364
rect 5037 10308 5093 10364
rect 5093 10308 5097 10364
rect 5033 10304 5097 10308
rect 5113 10364 5177 10368
rect 5113 10308 5117 10364
rect 5117 10308 5173 10364
rect 5173 10308 5177 10364
rect 5113 10304 5177 10308
rect 12715 10364 12779 10368
rect 12715 10308 12719 10364
rect 12719 10308 12775 10364
rect 12775 10308 12779 10364
rect 12715 10304 12779 10308
rect 12795 10364 12859 10368
rect 12795 10308 12799 10364
rect 12799 10308 12855 10364
rect 12855 10308 12859 10364
rect 12795 10304 12859 10308
rect 12875 10364 12939 10368
rect 12875 10308 12879 10364
rect 12879 10308 12935 10364
rect 12935 10308 12939 10364
rect 12875 10304 12939 10308
rect 12955 10364 13019 10368
rect 12955 10308 12959 10364
rect 12959 10308 13015 10364
rect 13015 10308 13019 10364
rect 12955 10304 13019 10308
rect 20557 10364 20621 10368
rect 20557 10308 20561 10364
rect 20561 10308 20617 10364
rect 20617 10308 20621 10364
rect 20557 10304 20621 10308
rect 20637 10364 20701 10368
rect 20637 10308 20641 10364
rect 20641 10308 20697 10364
rect 20697 10308 20701 10364
rect 20637 10304 20701 10308
rect 20717 10364 20781 10368
rect 20717 10308 20721 10364
rect 20721 10308 20777 10364
rect 20777 10308 20781 10364
rect 20717 10304 20781 10308
rect 20797 10364 20861 10368
rect 20797 10308 20801 10364
rect 20801 10308 20857 10364
rect 20857 10308 20861 10364
rect 20797 10304 20861 10308
rect 28399 10364 28463 10368
rect 28399 10308 28403 10364
rect 28403 10308 28459 10364
rect 28459 10308 28463 10364
rect 28399 10304 28463 10308
rect 28479 10364 28543 10368
rect 28479 10308 28483 10364
rect 28483 10308 28539 10364
rect 28539 10308 28543 10364
rect 28479 10304 28543 10308
rect 28559 10364 28623 10368
rect 28559 10308 28563 10364
rect 28563 10308 28619 10364
rect 28619 10308 28623 10364
rect 28559 10304 28623 10308
rect 28639 10364 28703 10368
rect 28639 10308 28643 10364
rect 28643 10308 28699 10364
rect 28699 10308 28703 10364
rect 28639 10304 28703 10308
rect 8794 9820 8858 9824
rect 8794 9764 8798 9820
rect 8798 9764 8854 9820
rect 8854 9764 8858 9820
rect 8794 9760 8858 9764
rect 8874 9820 8938 9824
rect 8874 9764 8878 9820
rect 8878 9764 8934 9820
rect 8934 9764 8938 9820
rect 8874 9760 8938 9764
rect 8954 9820 9018 9824
rect 8954 9764 8958 9820
rect 8958 9764 9014 9820
rect 9014 9764 9018 9820
rect 8954 9760 9018 9764
rect 9034 9820 9098 9824
rect 9034 9764 9038 9820
rect 9038 9764 9094 9820
rect 9094 9764 9098 9820
rect 9034 9760 9098 9764
rect 16636 9820 16700 9824
rect 16636 9764 16640 9820
rect 16640 9764 16696 9820
rect 16696 9764 16700 9820
rect 16636 9760 16700 9764
rect 16716 9820 16780 9824
rect 16716 9764 16720 9820
rect 16720 9764 16776 9820
rect 16776 9764 16780 9820
rect 16716 9760 16780 9764
rect 16796 9820 16860 9824
rect 16796 9764 16800 9820
rect 16800 9764 16856 9820
rect 16856 9764 16860 9820
rect 16796 9760 16860 9764
rect 16876 9820 16940 9824
rect 16876 9764 16880 9820
rect 16880 9764 16936 9820
rect 16936 9764 16940 9820
rect 16876 9760 16940 9764
rect 24478 9820 24542 9824
rect 24478 9764 24482 9820
rect 24482 9764 24538 9820
rect 24538 9764 24542 9820
rect 24478 9760 24542 9764
rect 24558 9820 24622 9824
rect 24558 9764 24562 9820
rect 24562 9764 24618 9820
rect 24618 9764 24622 9820
rect 24558 9760 24622 9764
rect 24638 9820 24702 9824
rect 24638 9764 24642 9820
rect 24642 9764 24698 9820
rect 24698 9764 24702 9820
rect 24638 9760 24702 9764
rect 24718 9820 24782 9824
rect 24718 9764 24722 9820
rect 24722 9764 24778 9820
rect 24778 9764 24782 9820
rect 24718 9760 24782 9764
rect 32320 9820 32384 9824
rect 32320 9764 32324 9820
rect 32324 9764 32380 9820
rect 32380 9764 32384 9820
rect 32320 9760 32384 9764
rect 32400 9820 32464 9824
rect 32400 9764 32404 9820
rect 32404 9764 32460 9820
rect 32460 9764 32464 9820
rect 32400 9760 32464 9764
rect 32480 9820 32544 9824
rect 32480 9764 32484 9820
rect 32484 9764 32540 9820
rect 32540 9764 32544 9820
rect 32480 9760 32544 9764
rect 32560 9820 32624 9824
rect 32560 9764 32564 9820
rect 32564 9764 32620 9820
rect 32620 9764 32624 9820
rect 32560 9760 32624 9764
rect 4873 9276 4937 9280
rect 4873 9220 4877 9276
rect 4877 9220 4933 9276
rect 4933 9220 4937 9276
rect 4873 9216 4937 9220
rect 4953 9276 5017 9280
rect 4953 9220 4957 9276
rect 4957 9220 5013 9276
rect 5013 9220 5017 9276
rect 4953 9216 5017 9220
rect 5033 9276 5097 9280
rect 5033 9220 5037 9276
rect 5037 9220 5093 9276
rect 5093 9220 5097 9276
rect 5033 9216 5097 9220
rect 5113 9276 5177 9280
rect 5113 9220 5117 9276
rect 5117 9220 5173 9276
rect 5173 9220 5177 9276
rect 5113 9216 5177 9220
rect 12715 9276 12779 9280
rect 12715 9220 12719 9276
rect 12719 9220 12775 9276
rect 12775 9220 12779 9276
rect 12715 9216 12779 9220
rect 12795 9276 12859 9280
rect 12795 9220 12799 9276
rect 12799 9220 12855 9276
rect 12855 9220 12859 9276
rect 12795 9216 12859 9220
rect 12875 9276 12939 9280
rect 12875 9220 12879 9276
rect 12879 9220 12935 9276
rect 12935 9220 12939 9276
rect 12875 9216 12939 9220
rect 12955 9276 13019 9280
rect 12955 9220 12959 9276
rect 12959 9220 13015 9276
rect 13015 9220 13019 9276
rect 12955 9216 13019 9220
rect 20557 9276 20621 9280
rect 20557 9220 20561 9276
rect 20561 9220 20617 9276
rect 20617 9220 20621 9276
rect 20557 9216 20621 9220
rect 20637 9276 20701 9280
rect 20637 9220 20641 9276
rect 20641 9220 20697 9276
rect 20697 9220 20701 9276
rect 20637 9216 20701 9220
rect 20717 9276 20781 9280
rect 20717 9220 20721 9276
rect 20721 9220 20777 9276
rect 20777 9220 20781 9276
rect 20717 9216 20781 9220
rect 20797 9276 20861 9280
rect 20797 9220 20801 9276
rect 20801 9220 20857 9276
rect 20857 9220 20861 9276
rect 20797 9216 20861 9220
rect 28399 9276 28463 9280
rect 28399 9220 28403 9276
rect 28403 9220 28459 9276
rect 28459 9220 28463 9276
rect 28399 9216 28463 9220
rect 28479 9276 28543 9280
rect 28479 9220 28483 9276
rect 28483 9220 28539 9276
rect 28539 9220 28543 9276
rect 28479 9216 28543 9220
rect 28559 9276 28623 9280
rect 28559 9220 28563 9276
rect 28563 9220 28619 9276
rect 28619 9220 28623 9276
rect 28559 9216 28623 9220
rect 28639 9276 28703 9280
rect 28639 9220 28643 9276
rect 28643 9220 28699 9276
rect 28699 9220 28703 9276
rect 28639 9216 28703 9220
rect 8794 8732 8858 8736
rect 8794 8676 8798 8732
rect 8798 8676 8854 8732
rect 8854 8676 8858 8732
rect 8794 8672 8858 8676
rect 8874 8732 8938 8736
rect 8874 8676 8878 8732
rect 8878 8676 8934 8732
rect 8934 8676 8938 8732
rect 8874 8672 8938 8676
rect 8954 8732 9018 8736
rect 8954 8676 8958 8732
rect 8958 8676 9014 8732
rect 9014 8676 9018 8732
rect 8954 8672 9018 8676
rect 9034 8732 9098 8736
rect 9034 8676 9038 8732
rect 9038 8676 9094 8732
rect 9094 8676 9098 8732
rect 9034 8672 9098 8676
rect 16636 8732 16700 8736
rect 16636 8676 16640 8732
rect 16640 8676 16696 8732
rect 16696 8676 16700 8732
rect 16636 8672 16700 8676
rect 16716 8732 16780 8736
rect 16716 8676 16720 8732
rect 16720 8676 16776 8732
rect 16776 8676 16780 8732
rect 16716 8672 16780 8676
rect 16796 8732 16860 8736
rect 16796 8676 16800 8732
rect 16800 8676 16856 8732
rect 16856 8676 16860 8732
rect 16796 8672 16860 8676
rect 16876 8732 16940 8736
rect 16876 8676 16880 8732
rect 16880 8676 16936 8732
rect 16936 8676 16940 8732
rect 16876 8672 16940 8676
rect 24478 8732 24542 8736
rect 24478 8676 24482 8732
rect 24482 8676 24538 8732
rect 24538 8676 24542 8732
rect 24478 8672 24542 8676
rect 24558 8732 24622 8736
rect 24558 8676 24562 8732
rect 24562 8676 24618 8732
rect 24618 8676 24622 8732
rect 24558 8672 24622 8676
rect 24638 8732 24702 8736
rect 24638 8676 24642 8732
rect 24642 8676 24698 8732
rect 24698 8676 24702 8732
rect 24638 8672 24702 8676
rect 24718 8732 24782 8736
rect 24718 8676 24722 8732
rect 24722 8676 24778 8732
rect 24778 8676 24782 8732
rect 24718 8672 24782 8676
rect 32320 8732 32384 8736
rect 32320 8676 32324 8732
rect 32324 8676 32380 8732
rect 32380 8676 32384 8732
rect 32320 8672 32384 8676
rect 32400 8732 32464 8736
rect 32400 8676 32404 8732
rect 32404 8676 32460 8732
rect 32460 8676 32464 8732
rect 32400 8672 32464 8676
rect 32480 8732 32544 8736
rect 32480 8676 32484 8732
rect 32484 8676 32540 8732
rect 32540 8676 32544 8732
rect 32480 8672 32544 8676
rect 32560 8732 32624 8736
rect 32560 8676 32564 8732
rect 32564 8676 32620 8732
rect 32620 8676 32624 8732
rect 32560 8672 32624 8676
rect 4873 8188 4937 8192
rect 4873 8132 4877 8188
rect 4877 8132 4933 8188
rect 4933 8132 4937 8188
rect 4873 8128 4937 8132
rect 4953 8188 5017 8192
rect 4953 8132 4957 8188
rect 4957 8132 5013 8188
rect 5013 8132 5017 8188
rect 4953 8128 5017 8132
rect 5033 8188 5097 8192
rect 5033 8132 5037 8188
rect 5037 8132 5093 8188
rect 5093 8132 5097 8188
rect 5033 8128 5097 8132
rect 5113 8188 5177 8192
rect 5113 8132 5117 8188
rect 5117 8132 5173 8188
rect 5173 8132 5177 8188
rect 5113 8128 5177 8132
rect 12715 8188 12779 8192
rect 12715 8132 12719 8188
rect 12719 8132 12775 8188
rect 12775 8132 12779 8188
rect 12715 8128 12779 8132
rect 12795 8188 12859 8192
rect 12795 8132 12799 8188
rect 12799 8132 12855 8188
rect 12855 8132 12859 8188
rect 12795 8128 12859 8132
rect 12875 8188 12939 8192
rect 12875 8132 12879 8188
rect 12879 8132 12935 8188
rect 12935 8132 12939 8188
rect 12875 8128 12939 8132
rect 12955 8188 13019 8192
rect 12955 8132 12959 8188
rect 12959 8132 13015 8188
rect 13015 8132 13019 8188
rect 12955 8128 13019 8132
rect 20557 8188 20621 8192
rect 20557 8132 20561 8188
rect 20561 8132 20617 8188
rect 20617 8132 20621 8188
rect 20557 8128 20621 8132
rect 20637 8188 20701 8192
rect 20637 8132 20641 8188
rect 20641 8132 20697 8188
rect 20697 8132 20701 8188
rect 20637 8128 20701 8132
rect 20717 8188 20781 8192
rect 20717 8132 20721 8188
rect 20721 8132 20777 8188
rect 20777 8132 20781 8188
rect 20717 8128 20781 8132
rect 20797 8188 20861 8192
rect 20797 8132 20801 8188
rect 20801 8132 20857 8188
rect 20857 8132 20861 8188
rect 20797 8128 20861 8132
rect 28399 8188 28463 8192
rect 28399 8132 28403 8188
rect 28403 8132 28459 8188
rect 28459 8132 28463 8188
rect 28399 8128 28463 8132
rect 28479 8188 28543 8192
rect 28479 8132 28483 8188
rect 28483 8132 28539 8188
rect 28539 8132 28543 8188
rect 28479 8128 28543 8132
rect 28559 8188 28623 8192
rect 28559 8132 28563 8188
rect 28563 8132 28619 8188
rect 28619 8132 28623 8188
rect 28559 8128 28623 8132
rect 28639 8188 28703 8192
rect 28639 8132 28643 8188
rect 28643 8132 28699 8188
rect 28699 8132 28703 8188
rect 28639 8128 28703 8132
rect 8794 7644 8858 7648
rect 8794 7588 8798 7644
rect 8798 7588 8854 7644
rect 8854 7588 8858 7644
rect 8794 7584 8858 7588
rect 8874 7644 8938 7648
rect 8874 7588 8878 7644
rect 8878 7588 8934 7644
rect 8934 7588 8938 7644
rect 8874 7584 8938 7588
rect 8954 7644 9018 7648
rect 8954 7588 8958 7644
rect 8958 7588 9014 7644
rect 9014 7588 9018 7644
rect 8954 7584 9018 7588
rect 9034 7644 9098 7648
rect 9034 7588 9038 7644
rect 9038 7588 9094 7644
rect 9094 7588 9098 7644
rect 9034 7584 9098 7588
rect 16636 7644 16700 7648
rect 16636 7588 16640 7644
rect 16640 7588 16696 7644
rect 16696 7588 16700 7644
rect 16636 7584 16700 7588
rect 16716 7644 16780 7648
rect 16716 7588 16720 7644
rect 16720 7588 16776 7644
rect 16776 7588 16780 7644
rect 16716 7584 16780 7588
rect 16796 7644 16860 7648
rect 16796 7588 16800 7644
rect 16800 7588 16856 7644
rect 16856 7588 16860 7644
rect 16796 7584 16860 7588
rect 16876 7644 16940 7648
rect 16876 7588 16880 7644
rect 16880 7588 16936 7644
rect 16936 7588 16940 7644
rect 16876 7584 16940 7588
rect 24478 7644 24542 7648
rect 24478 7588 24482 7644
rect 24482 7588 24538 7644
rect 24538 7588 24542 7644
rect 24478 7584 24542 7588
rect 24558 7644 24622 7648
rect 24558 7588 24562 7644
rect 24562 7588 24618 7644
rect 24618 7588 24622 7644
rect 24558 7584 24622 7588
rect 24638 7644 24702 7648
rect 24638 7588 24642 7644
rect 24642 7588 24698 7644
rect 24698 7588 24702 7644
rect 24638 7584 24702 7588
rect 24718 7644 24782 7648
rect 24718 7588 24722 7644
rect 24722 7588 24778 7644
rect 24778 7588 24782 7644
rect 24718 7584 24782 7588
rect 32320 7644 32384 7648
rect 32320 7588 32324 7644
rect 32324 7588 32380 7644
rect 32380 7588 32384 7644
rect 32320 7584 32384 7588
rect 32400 7644 32464 7648
rect 32400 7588 32404 7644
rect 32404 7588 32460 7644
rect 32460 7588 32464 7644
rect 32400 7584 32464 7588
rect 32480 7644 32544 7648
rect 32480 7588 32484 7644
rect 32484 7588 32540 7644
rect 32540 7588 32544 7644
rect 32480 7584 32544 7588
rect 32560 7644 32624 7648
rect 32560 7588 32564 7644
rect 32564 7588 32620 7644
rect 32620 7588 32624 7644
rect 32560 7584 32624 7588
rect 4873 7100 4937 7104
rect 4873 7044 4877 7100
rect 4877 7044 4933 7100
rect 4933 7044 4937 7100
rect 4873 7040 4937 7044
rect 4953 7100 5017 7104
rect 4953 7044 4957 7100
rect 4957 7044 5013 7100
rect 5013 7044 5017 7100
rect 4953 7040 5017 7044
rect 5033 7100 5097 7104
rect 5033 7044 5037 7100
rect 5037 7044 5093 7100
rect 5093 7044 5097 7100
rect 5033 7040 5097 7044
rect 5113 7100 5177 7104
rect 5113 7044 5117 7100
rect 5117 7044 5173 7100
rect 5173 7044 5177 7100
rect 5113 7040 5177 7044
rect 12715 7100 12779 7104
rect 12715 7044 12719 7100
rect 12719 7044 12775 7100
rect 12775 7044 12779 7100
rect 12715 7040 12779 7044
rect 12795 7100 12859 7104
rect 12795 7044 12799 7100
rect 12799 7044 12855 7100
rect 12855 7044 12859 7100
rect 12795 7040 12859 7044
rect 12875 7100 12939 7104
rect 12875 7044 12879 7100
rect 12879 7044 12935 7100
rect 12935 7044 12939 7100
rect 12875 7040 12939 7044
rect 12955 7100 13019 7104
rect 12955 7044 12959 7100
rect 12959 7044 13015 7100
rect 13015 7044 13019 7100
rect 12955 7040 13019 7044
rect 20557 7100 20621 7104
rect 20557 7044 20561 7100
rect 20561 7044 20617 7100
rect 20617 7044 20621 7100
rect 20557 7040 20621 7044
rect 20637 7100 20701 7104
rect 20637 7044 20641 7100
rect 20641 7044 20697 7100
rect 20697 7044 20701 7100
rect 20637 7040 20701 7044
rect 20717 7100 20781 7104
rect 20717 7044 20721 7100
rect 20721 7044 20777 7100
rect 20777 7044 20781 7100
rect 20717 7040 20781 7044
rect 20797 7100 20861 7104
rect 20797 7044 20801 7100
rect 20801 7044 20857 7100
rect 20857 7044 20861 7100
rect 20797 7040 20861 7044
rect 28399 7100 28463 7104
rect 28399 7044 28403 7100
rect 28403 7044 28459 7100
rect 28459 7044 28463 7100
rect 28399 7040 28463 7044
rect 28479 7100 28543 7104
rect 28479 7044 28483 7100
rect 28483 7044 28539 7100
rect 28539 7044 28543 7100
rect 28479 7040 28543 7044
rect 28559 7100 28623 7104
rect 28559 7044 28563 7100
rect 28563 7044 28619 7100
rect 28619 7044 28623 7100
rect 28559 7040 28623 7044
rect 28639 7100 28703 7104
rect 28639 7044 28643 7100
rect 28643 7044 28699 7100
rect 28699 7044 28703 7100
rect 28639 7040 28703 7044
rect 8794 6556 8858 6560
rect 8794 6500 8798 6556
rect 8798 6500 8854 6556
rect 8854 6500 8858 6556
rect 8794 6496 8858 6500
rect 8874 6556 8938 6560
rect 8874 6500 8878 6556
rect 8878 6500 8934 6556
rect 8934 6500 8938 6556
rect 8874 6496 8938 6500
rect 8954 6556 9018 6560
rect 8954 6500 8958 6556
rect 8958 6500 9014 6556
rect 9014 6500 9018 6556
rect 8954 6496 9018 6500
rect 9034 6556 9098 6560
rect 9034 6500 9038 6556
rect 9038 6500 9094 6556
rect 9094 6500 9098 6556
rect 9034 6496 9098 6500
rect 16636 6556 16700 6560
rect 16636 6500 16640 6556
rect 16640 6500 16696 6556
rect 16696 6500 16700 6556
rect 16636 6496 16700 6500
rect 16716 6556 16780 6560
rect 16716 6500 16720 6556
rect 16720 6500 16776 6556
rect 16776 6500 16780 6556
rect 16716 6496 16780 6500
rect 16796 6556 16860 6560
rect 16796 6500 16800 6556
rect 16800 6500 16856 6556
rect 16856 6500 16860 6556
rect 16796 6496 16860 6500
rect 16876 6556 16940 6560
rect 16876 6500 16880 6556
rect 16880 6500 16936 6556
rect 16936 6500 16940 6556
rect 16876 6496 16940 6500
rect 24478 6556 24542 6560
rect 24478 6500 24482 6556
rect 24482 6500 24538 6556
rect 24538 6500 24542 6556
rect 24478 6496 24542 6500
rect 24558 6556 24622 6560
rect 24558 6500 24562 6556
rect 24562 6500 24618 6556
rect 24618 6500 24622 6556
rect 24558 6496 24622 6500
rect 24638 6556 24702 6560
rect 24638 6500 24642 6556
rect 24642 6500 24698 6556
rect 24698 6500 24702 6556
rect 24638 6496 24702 6500
rect 24718 6556 24782 6560
rect 24718 6500 24722 6556
rect 24722 6500 24778 6556
rect 24778 6500 24782 6556
rect 24718 6496 24782 6500
rect 32320 6556 32384 6560
rect 32320 6500 32324 6556
rect 32324 6500 32380 6556
rect 32380 6500 32384 6556
rect 32320 6496 32384 6500
rect 32400 6556 32464 6560
rect 32400 6500 32404 6556
rect 32404 6500 32460 6556
rect 32460 6500 32464 6556
rect 32400 6496 32464 6500
rect 32480 6556 32544 6560
rect 32480 6500 32484 6556
rect 32484 6500 32540 6556
rect 32540 6500 32544 6556
rect 32480 6496 32544 6500
rect 32560 6556 32624 6560
rect 32560 6500 32564 6556
rect 32564 6500 32620 6556
rect 32620 6500 32624 6556
rect 32560 6496 32624 6500
rect 4873 6012 4937 6016
rect 4873 5956 4877 6012
rect 4877 5956 4933 6012
rect 4933 5956 4937 6012
rect 4873 5952 4937 5956
rect 4953 6012 5017 6016
rect 4953 5956 4957 6012
rect 4957 5956 5013 6012
rect 5013 5956 5017 6012
rect 4953 5952 5017 5956
rect 5033 6012 5097 6016
rect 5033 5956 5037 6012
rect 5037 5956 5093 6012
rect 5093 5956 5097 6012
rect 5033 5952 5097 5956
rect 5113 6012 5177 6016
rect 5113 5956 5117 6012
rect 5117 5956 5173 6012
rect 5173 5956 5177 6012
rect 5113 5952 5177 5956
rect 12715 6012 12779 6016
rect 12715 5956 12719 6012
rect 12719 5956 12775 6012
rect 12775 5956 12779 6012
rect 12715 5952 12779 5956
rect 12795 6012 12859 6016
rect 12795 5956 12799 6012
rect 12799 5956 12855 6012
rect 12855 5956 12859 6012
rect 12795 5952 12859 5956
rect 12875 6012 12939 6016
rect 12875 5956 12879 6012
rect 12879 5956 12935 6012
rect 12935 5956 12939 6012
rect 12875 5952 12939 5956
rect 12955 6012 13019 6016
rect 12955 5956 12959 6012
rect 12959 5956 13015 6012
rect 13015 5956 13019 6012
rect 12955 5952 13019 5956
rect 20557 6012 20621 6016
rect 20557 5956 20561 6012
rect 20561 5956 20617 6012
rect 20617 5956 20621 6012
rect 20557 5952 20621 5956
rect 20637 6012 20701 6016
rect 20637 5956 20641 6012
rect 20641 5956 20697 6012
rect 20697 5956 20701 6012
rect 20637 5952 20701 5956
rect 20717 6012 20781 6016
rect 20717 5956 20721 6012
rect 20721 5956 20777 6012
rect 20777 5956 20781 6012
rect 20717 5952 20781 5956
rect 20797 6012 20861 6016
rect 20797 5956 20801 6012
rect 20801 5956 20857 6012
rect 20857 5956 20861 6012
rect 20797 5952 20861 5956
rect 28399 6012 28463 6016
rect 28399 5956 28403 6012
rect 28403 5956 28459 6012
rect 28459 5956 28463 6012
rect 28399 5952 28463 5956
rect 28479 6012 28543 6016
rect 28479 5956 28483 6012
rect 28483 5956 28539 6012
rect 28539 5956 28543 6012
rect 28479 5952 28543 5956
rect 28559 6012 28623 6016
rect 28559 5956 28563 6012
rect 28563 5956 28619 6012
rect 28619 5956 28623 6012
rect 28559 5952 28623 5956
rect 28639 6012 28703 6016
rect 28639 5956 28643 6012
rect 28643 5956 28699 6012
rect 28699 5956 28703 6012
rect 28639 5952 28703 5956
rect 8794 5468 8858 5472
rect 8794 5412 8798 5468
rect 8798 5412 8854 5468
rect 8854 5412 8858 5468
rect 8794 5408 8858 5412
rect 8874 5468 8938 5472
rect 8874 5412 8878 5468
rect 8878 5412 8934 5468
rect 8934 5412 8938 5468
rect 8874 5408 8938 5412
rect 8954 5468 9018 5472
rect 8954 5412 8958 5468
rect 8958 5412 9014 5468
rect 9014 5412 9018 5468
rect 8954 5408 9018 5412
rect 9034 5468 9098 5472
rect 9034 5412 9038 5468
rect 9038 5412 9094 5468
rect 9094 5412 9098 5468
rect 9034 5408 9098 5412
rect 16636 5468 16700 5472
rect 16636 5412 16640 5468
rect 16640 5412 16696 5468
rect 16696 5412 16700 5468
rect 16636 5408 16700 5412
rect 16716 5468 16780 5472
rect 16716 5412 16720 5468
rect 16720 5412 16776 5468
rect 16776 5412 16780 5468
rect 16716 5408 16780 5412
rect 16796 5468 16860 5472
rect 16796 5412 16800 5468
rect 16800 5412 16856 5468
rect 16856 5412 16860 5468
rect 16796 5408 16860 5412
rect 16876 5468 16940 5472
rect 16876 5412 16880 5468
rect 16880 5412 16936 5468
rect 16936 5412 16940 5468
rect 16876 5408 16940 5412
rect 24478 5468 24542 5472
rect 24478 5412 24482 5468
rect 24482 5412 24538 5468
rect 24538 5412 24542 5468
rect 24478 5408 24542 5412
rect 24558 5468 24622 5472
rect 24558 5412 24562 5468
rect 24562 5412 24618 5468
rect 24618 5412 24622 5468
rect 24558 5408 24622 5412
rect 24638 5468 24702 5472
rect 24638 5412 24642 5468
rect 24642 5412 24698 5468
rect 24698 5412 24702 5468
rect 24638 5408 24702 5412
rect 24718 5468 24782 5472
rect 24718 5412 24722 5468
rect 24722 5412 24778 5468
rect 24778 5412 24782 5468
rect 24718 5408 24782 5412
rect 32320 5468 32384 5472
rect 32320 5412 32324 5468
rect 32324 5412 32380 5468
rect 32380 5412 32384 5468
rect 32320 5408 32384 5412
rect 32400 5468 32464 5472
rect 32400 5412 32404 5468
rect 32404 5412 32460 5468
rect 32460 5412 32464 5468
rect 32400 5408 32464 5412
rect 32480 5468 32544 5472
rect 32480 5412 32484 5468
rect 32484 5412 32540 5468
rect 32540 5412 32544 5468
rect 32480 5408 32544 5412
rect 32560 5468 32624 5472
rect 32560 5412 32564 5468
rect 32564 5412 32620 5468
rect 32620 5412 32624 5468
rect 32560 5408 32624 5412
rect 4873 4924 4937 4928
rect 4873 4868 4877 4924
rect 4877 4868 4933 4924
rect 4933 4868 4937 4924
rect 4873 4864 4937 4868
rect 4953 4924 5017 4928
rect 4953 4868 4957 4924
rect 4957 4868 5013 4924
rect 5013 4868 5017 4924
rect 4953 4864 5017 4868
rect 5033 4924 5097 4928
rect 5033 4868 5037 4924
rect 5037 4868 5093 4924
rect 5093 4868 5097 4924
rect 5033 4864 5097 4868
rect 5113 4924 5177 4928
rect 5113 4868 5117 4924
rect 5117 4868 5173 4924
rect 5173 4868 5177 4924
rect 5113 4864 5177 4868
rect 12715 4924 12779 4928
rect 12715 4868 12719 4924
rect 12719 4868 12775 4924
rect 12775 4868 12779 4924
rect 12715 4864 12779 4868
rect 12795 4924 12859 4928
rect 12795 4868 12799 4924
rect 12799 4868 12855 4924
rect 12855 4868 12859 4924
rect 12795 4864 12859 4868
rect 12875 4924 12939 4928
rect 12875 4868 12879 4924
rect 12879 4868 12935 4924
rect 12935 4868 12939 4924
rect 12875 4864 12939 4868
rect 12955 4924 13019 4928
rect 12955 4868 12959 4924
rect 12959 4868 13015 4924
rect 13015 4868 13019 4924
rect 12955 4864 13019 4868
rect 20557 4924 20621 4928
rect 20557 4868 20561 4924
rect 20561 4868 20617 4924
rect 20617 4868 20621 4924
rect 20557 4864 20621 4868
rect 20637 4924 20701 4928
rect 20637 4868 20641 4924
rect 20641 4868 20697 4924
rect 20697 4868 20701 4924
rect 20637 4864 20701 4868
rect 20717 4924 20781 4928
rect 20717 4868 20721 4924
rect 20721 4868 20777 4924
rect 20777 4868 20781 4924
rect 20717 4864 20781 4868
rect 20797 4924 20861 4928
rect 20797 4868 20801 4924
rect 20801 4868 20857 4924
rect 20857 4868 20861 4924
rect 20797 4864 20861 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 28639 4924 28703 4928
rect 28639 4868 28643 4924
rect 28643 4868 28699 4924
rect 28699 4868 28703 4924
rect 28639 4864 28703 4868
rect 8794 4380 8858 4384
rect 8794 4324 8798 4380
rect 8798 4324 8854 4380
rect 8854 4324 8858 4380
rect 8794 4320 8858 4324
rect 8874 4380 8938 4384
rect 8874 4324 8878 4380
rect 8878 4324 8934 4380
rect 8934 4324 8938 4380
rect 8874 4320 8938 4324
rect 8954 4380 9018 4384
rect 8954 4324 8958 4380
rect 8958 4324 9014 4380
rect 9014 4324 9018 4380
rect 8954 4320 9018 4324
rect 9034 4380 9098 4384
rect 9034 4324 9038 4380
rect 9038 4324 9094 4380
rect 9094 4324 9098 4380
rect 9034 4320 9098 4324
rect 16636 4380 16700 4384
rect 16636 4324 16640 4380
rect 16640 4324 16696 4380
rect 16696 4324 16700 4380
rect 16636 4320 16700 4324
rect 16716 4380 16780 4384
rect 16716 4324 16720 4380
rect 16720 4324 16776 4380
rect 16776 4324 16780 4380
rect 16716 4320 16780 4324
rect 16796 4380 16860 4384
rect 16796 4324 16800 4380
rect 16800 4324 16856 4380
rect 16856 4324 16860 4380
rect 16796 4320 16860 4324
rect 16876 4380 16940 4384
rect 16876 4324 16880 4380
rect 16880 4324 16936 4380
rect 16936 4324 16940 4380
rect 16876 4320 16940 4324
rect 24478 4380 24542 4384
rect 24478 4324 24482 4380
rect 24482 4324 24538 4380
rect 24538 4324 24542 4380
rect 24478 4320 24542 4324
rect 24558 4380 24622 4384
rect 24558 4324 24562 4380
rect 24562 4324 24618 4380
rect 24618 4324 24622 4380
rect 24558 4320 24622 4324
rect 24638 4380 24702 4384
rect 24638 4324 24642 4380
rect 24642 4324 24698 4380
rect 24698 4324 24702 4380
rect 24638 4320 24702 4324
rect 24718 4380 24782 4384
rect 24718 4324 24722 4380
rect 24722 4324 24778 4380
rect 24778 4324 24782 4380
rect 24718 4320 24782 4324
rect 32320 4380 32384 4384
rect 32320 4324 32324 4380
rect 32324 4324 32380 4380
rect 32380 4324 32384 4380
rect 32320 4320 32384 4324
rect 32400 4380 32464 4384
rect 32400 4324 32404 4380
rect 32404 4324 32460 4380
rect 32460 4324 32464 4380
rect 32400 4320 32464 4324
rect 32480 4380 32544 4384
rect 32480 4324 32484 4380
rect 32484 4324 32540 4380
rect 32540 4324 32544 4380
rect 32480 4320 32544 4324
rect 32560 4380 32624 4384
rect 32560 4324 32564 4380
rect 32564 4324 32620 4380
rect 32620 4324 32624 4380
rect 32560 4320 32624 4324
rect 4873 3836 4937 3840
rect 4873 3780 4877 3836
rect 4877 3780 4933 3836
rect 4933 3780 4937 3836
rect 4873 3776 4937 3780
rect 4953 3836 5017 3840
rect 4953 3780 4957 3836
rect 4957 3780 5013 3836
rect 5013 3780 5017 3836
rect 4953 3776 5017 3780
rect 5033 3836 5097 3840
rect 5033 3780 5037 3836
rect 5037 3780 5093 3836
rect 5093 3780 5097 3836
rect 5033 3776 5097 3780
rect 5113 3836 5177 3840
rect 5113 3780 5117 3836
rect 5117 3780 5173 3836
rect 5173 3780 5177 3836
rect 5113 3776 5177 3780
rect 12715 3836 12779 3840
rect 12715 3780 12719 3836
rect 12719 3780 12775 3836
rect 12775 3780 12779 3836
rect 12715 3776 12779 3780
rect 12795 3836 12859 3840
rect 12795 3780 12799 3836
rect 12799 3780 12855 3836
rect 12855 3780 12859 3836
rect 12795 3776 12859 3780
rect 12875 3836 12939 3840
rect 12875 3780 12879 3836
rect 12879 3780 12935 3836
rect 12935 3780 12939 3836
rect 12875 3776 12939 3780
rect 12955 3836 13019 3840
rect 12955 3780 12959 3836
rect 12959 3780 13015 3836
rect 13015 3780 13019 3836
rect 12955 3776 13019 3780
rect 20557 3836 20621 3840
rect 20557 3780 20561 3836
rect 20561 3780 20617 3836
rect 20617 3780 20621 3836
rect 20557 3776 20621 3780
rect 20637 3836 20701 3840
rect 20637 3780 20641 3836
rect 20641 3780 20697 3836
rect 20697 3780 20701 3836
rect 20637 3776 20701 3780
rect 20717 3836 20781 3840
rect 20717 3780 20721 3836
rect 20721 3780 20777 3836
rect 20777 3780 20781 3836
rect 20717 3776 20781 3780
rect 20797 3836 20861 3840
rect 20797 3780 20801 3836
rect 20801 3780 20857 3836
rect 20857 3780 20861 3836
rect 20797 3776 20861 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 28639 3836 28703 3840
rect 28639 3780 28643 3836
rect 28643 3780 28699 3836
rect 28699 3780 28703 3836
rect 28639 3776 28703 3780
rect 8794 3292 8858 3296
rect 8794 3236 8798 3292
rect 8798 3236 8854 3292
rect 8854 3236 8858 3292
rect 8794 3232 8858 3236
rect 8874 3292 8938 3296
rect 8874 3236 8878 3292
rect 8878 3236 8934 3292
rect 8934 3236 8938 3292
rect 8874 3232 8938 3236
rect 8954 3292 9018 3296
rect 8954 3236 8958 3292
rect 8958 3236 9014 3292
rect 9014 3236 9018 3292
rect 8954 3232 9018 3236
rect 9034 3292 9098 3296
rect 9034 3236 9038 3292
rect 9038 3236 9094 3292
rect 9094 3236 9098 3292
rect 9034 3232 9098 3236
rect 16636 3292 16700 3296
rect 16636 3236 16640 3292
rect 16640 3236 16696 3292
rect 16696 3236 16700 3292
rect 16636 3232 16700 3236
rect 16716 3292 16780 3296
rect 16716 3236 16720 3292
rect 16720 3236 16776 3292
rect 16776 3236 16780 3292
rect 16716 3232 16780 3236
rect 16796 3292 16860 3296
rect 16796 3236 16800 3292
rect 16800 3236 16856 3292
rect 16856 3236 16860 3292
rect 16796 3232 16860 3236
rect 16876 3292 16940 3296
rect 16876 3236 16880 3292
rect 16880 3236 16936 3292
rect 16936 3236 16940 3292
rect 16876 3232 16940 3236
rect 24478 3292 24542 3296
rect 24478 3236 24482 3292
rect 24482 3236 24538 3292
rect 24538 3236 24542 3292
rect 24478 3232 24542 3236
rect 24558 3292 24622 3296
rect 24558 3236 24562 3292
rect 24562 3236 24618 3292
rect 24618 3236 24622 3292
rect 24558 3232 24622 3236
rect 24638 3292 24702 3296
rect 24638 3236 24642 3292
rect 24642 3236 24698 3292
rect 24698 3236 24702 3292
rect 24638 3232 24702 3236
rect 24718 3292 24782 3296
rect 24718 3236 24722 3292
rect 24722 3236 24778 3292
rect 24778 3236 24782 3292
rect 24718 3232 24782 3236
rect 32320 3292 32384 3296
rect 32320 3236 32324 3292
rect 32324 3236 32380 3292
rect 32380 3236 32384 3292
rect 32320 3232 32384 3236
rect 32400 3292 32464 3296
rect 32400 3236 32404 3292
rect 32404 3236 32460 3292
rect 32460 3236 32464 3292
rect 32400 3232 32464 3236
rect 32480 3292 32544 3296
rect 32480 3236 32484 3292
rect 32484 3236 32540 3292
rect 32540 3236 32544 3292
rect 32480 3232 32544 3236
rect 32560 3292 32624 3296
rect 32560 3236 32564 3292
rect 32564 3236 32620 3292
rect 32620 3236 32624 3292
rect 32560 3232 32624 3236
rect 4873 2748 4937 2752
rect 4873 2692 4877 2748
rect 4877 2692 4933 2748
rect 4933 2692 4937 2748
rect 4873 2688 4937 2692
rect 4953 2748 5017 2752
rect 4953 2692 4957 2748
rect 4957 2692 5013 2748
rect 5013 2692 5017 2748
rect 4953 2688 5017 2692
rect 5033 2748 5097 2752
rect 5033 2692 5037 2748
rect 5037 2692 5093 2748
rect 5093 2692 5097 2748
rect 5033 2688 5097 2692
rect 5113 2748 5177 2752
rect 5113 2692 5117 2748
rect 5117 2692 5173 2748
rect 5173 2692 5177 2748
rect 5113 2688 5177 2692
rect 12715 2748 12779 2752
rect 12715 2692 12719 2748
rect 12719 2692 12775 2748
rect 12775 2692 12779 2748
rect 12715 2688 12779 2692
rect 12795 2748 12859 2752
rect 12795 2692 12799 2748
rect 12799 2692 12855 2748
rect 12855 2692 12859 2748
rect 12795 2688 12859 2692
rect 12875 2748 12939 2752
rect 12875 2692 12879 2748
rect 12879 2692 12935 2748
rect 12935 2692 12939 2748
rect 12875 2688 12939 2692
rect 12955 2748 13019 2752
rect 12955 2692 12959 2748
rect 12959 2692 13015 2748
rect 13015 2692 13019 2748
rect 12955 2688 13019 2692
rect 20557 2748 20621 2752
rect 20557 2692 20561 2748
rect 20561 2692 20617 2748
rect 20617 2692 20621 2748
rect 20557 2688 20621 2692
rect 20637 2748 20701 2752
rect 20637 2692 20641 2748
rect 20641 2692 20697 2748
rect 20697 2692 20701 2748
rect 20637 2688 20701 2692
rect 20717 2748 20781 2752
rect 20717 2692 20721 2748
rect 20721 2692 20777 2748
rect 20777 2692 20781 2748
rect 20717 2688 20781 2692
rect 20797 2748 20861 2752
rect 20797 2692 20801 2748
rect 20801 2692 20857 2748
rect 20857 2692 20861 2748
rect 20797 2688 20861 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 28639 2748 28703 2752
rect 28639 2692 28643 2748
rect 28643 2692 28699 2748
rect 28699 2692 28703 2748
rect 28639 2688 28703 2692
rect 8794 2204 8858 2208
rect 8794 2148 8798 2204
rect 8798 2148 8854 2204
rect 8854 2148 8858 2204
rect 8794 2144 8858 2148
rect 8874 2204 8938 2208
rect 8874 2148 8878 2204
rect 8878 2148 8934 2204
rect 8934 2148 8938 2204
rect 8874 2144 8938 2148
rect 8954 2204 9018 2208
rect 8954 2148 8958 2204
rect 8958 2148 9014 2204
rect 9014 2148 9018 2204
rect 8954 2144 9018 2148
rect 9034 2204 9098 2208
rect 9034 2148 9038 2204
rect 9038 2148 9094 2204
rect 9094 2148 9098 2204
rect 9034 2144 9098 2148
rect 16636 2204 16700 2208
rect 16636 2148 16640 2204
rect 16640 2148 16696 2204
rect 16696 2148 16700 2204
rect 16636 2144 16700 2148
rect 16716 2204 16780 2208
rect 16716 2148 16720 2204
rect 16720 2148 16776 2204
rect 16776 2148 16780 2204
rect 16716 2144 16780 2148
rect 16796 2204 16860 2208
rect 16796 2148 16800 2204
rect 16800 2148 16856 2204
rect 16856 2148 16860 2204
rect 16796 2144 16860 2148
rect 16876 2204 16940 2208
rect 16876 2148 16880 2204
rect 16880 2148 16936 2204
rect 16936 2148 16940 2204
rect 16876 2144 16940 2148
rect 24478 2204 24542 2208
rect 24478 2148 24482 2204
rect 24482 2148 24538 2204
rect 24538 2148 24542 2204
rect 24478 2144 24542 2148
rect 24558 2204 24622 2208
rect 24558 2148 24562 2204
rect 24562 2148 24618 2204
rect 24618 2148 24622 2204
rect 24558 2144 24622 2148
rect 24638 2204 24702 2208
rect 24638 2148 24642 2204
rect 24642 2148 24698 2204
rect 24698 2148 24702 2204
rect 24638 2144 24702 2148
rect 24718 2204 24782 2208
rect 24718 2148 24722 2204
rect 24722 2148 24778 2204
rect 24778 2148 24782 2204
rect 24718 2144 24782 2148
rect 32320 2204 32384 2208
rect 32320 2148 32324 2204
rect 32324 2148 32380 2204
rect 32380 2148 32384 2204
rect 32320 2144 32384 2148
rect 32400 2204 32464 2208
rect 32400 2148 32404 2204
rect 32404 2148 32460 2204
rect 32460 2148 32464 2204
rect 32400 2144 32464 2148
rect 32480 2204 32544 2208
rect 32480 2148 32484 2204
rect 32484 2148 32540 2204
rect 32540 2148 32544 2204
rect 32480 2144 32544 2148
rect 32560 2204 32624 2208
rect 32560 2148 32564 2204
rect 32564 2148 32620 2204
rect 32620 2148 32624 2204
rect 32560 2144 32624 2148
rect 4873 1660 4937 1664
rect 4873 1604 4877 1660
rect 4877 1604 4933 1660
rect 4933 1604 4937 1660
rect 4873 1600 4937 1604
rect 4953 1660 5017 1664
rect 4953 1604 4957 1660
rect 4957 1604 5013 1660
rect 5013 1604 5017 1660
rect 4953 1600 5017 1604
rect 5033 1660 5097 1664
rect 5033 1604 5037 1660
rect 5037 1604 5093 1660
rect 5093 1604 5097 1660
rect 5033 1600 5097 1604
rect 5113 1660 5177 1664
rect 5113 1604 5117 1660
rect 5117 1604 5173 1660
rect 5173 1604 5177 1660
rect 5113 1600 5177 1604
rect 12715 1660 12779 1664
rect 12715 1604 12719 1660
rect 12719 1604 12775 1660
rect 12775 1604 12779 1660
rect 12715 1600 12779 1604
rect 12795 1660 12859 1664
rect 12795 1604 12799 1660
rect 12799 1604 12855 1660
rect 12855 1604 12859 1660
rect 12795 1600 12859 1604
rect 12875 1660 12939 1664
rect 12875 1604 12879 1660
rect 12879 1604 12935 1660
rect 12935 1604 12939 1660
rect 12875 1600 12939 1604
rect 12955 1660 13019 1664
rect 12955 1604 12959 1660
rect 12959 1604 13015 1660
rect 13015 1604 13019 1660
rect 12955 1600 13019 1604
rect 20557 1660 20621 1664
rect 20557 1604 20561 1660
rect 20561 1604 20617 1660
rect 20617 1604 20621 1660
rect 20557 1600 20621 1604
rect 20637 1660 20701 1664
rect 20637 1604 20641 1660
rect 20641 1604 20697 1660
rect 20697 1604 20701 1660
rect 20637 1600 20701 1604
rect 20717 1660 20781 1664
rect 20717 1604 20721 1660
rect 20721 1604 20777 1660
rect 20777 1604 20781 1660
rect 20717 1600 20781 1604
rect 20797 1660 20861 1664
rect 20797 1604 20801 1660
rect 20801 1604 20857 1660
rect 20857 1604 20861 1660
rect 20797 1600 20861 1604
rect 28399 1660 28463 1664
rect 28399 1604 28403 1660
rect 28403 1604 28459 1660
rect 28459 1604 28463 1660
rect 28399 1600 28463 1604
rect 28479 1660 28543 1664
rect 28479 1604 28483 1660
rect 28483 1604 28539 1660
rect 28539 1604 28543 1660
rect 28479 1600 28543 1604
rect 28559 1660 28623 1664
rect 28559 1604 28563 1660
rect 28563 1604 28619 1660
rect 28619 1604 28623 1660
rect 28559 1600 28623 1604
rect 28639 1660 28703 1664
rect 28639 1604 28643 1660
rect 28643 1604 28699 1660
rect 28699 1604 28703 1660
rect 28639 1600 28703 1604
rect 8794 1116 8858 1120
rect 8794 1060 8798 1116
rect 8798 1060 8854 1116
rect 8854 1060 8858 1116
rect 8794 1056 8858 1060
rect 8874 1116 8938 1120
rect 8874 1060 8878 1116
rect 8878 1060 8934 1116
rect 8934 1060 8938 1116
rect 8874 1056 8938 1060
rect 8954 1116 9018 1120
rect 8954 1060 8958 1116
rect 8958 1060 9014 1116
rect 9014 1060 9018 1116
rect 8954 1056 9018 1060
rect 9034 1116 9098 1120
rect 9034 1060 9038 1116
rect 9038 1060 9094 1116
rect 9094 1060 9098 1116
rect 9034 1056 9098 1060
rect 16636 1116 16700 1120
rect 16636 1060 16640 1116
rect 16640 1060 16696 1116
rect 16696 1060 16700 1116
rect 16636 1056 16700 1060
rect 16716 1116 16780 1120
rect 16716 1060 16720 1116
rect 16720 1060 16776 1116
rect 16776 1060 16780 1116
rect 16716 1056 16780 1060
rect 16796 1116 16860 1120
rect 16796 1060 16800 1116
rect 16800 1060 16856 1116
rect 16856 1060 16860 1116
rect 16796 1056 16860 1060
rect 16876 1116 16940 1120
rect 16876 1060 16880 1116
rect 16880 1060 16936 1116
rect 16936 1060 16940 1116
rect 16876 1056 16940 1060
rect 24478 1116 24542 1120
rect 24478 1060 24482 1116
rect 24482 1060 24538 1116
rect 24538 1060 24542 1116
rect 24478 1056 24542 1060
rect 24558 1116 24622 1120
rect 24558 1060 24562 1116
rect 24562 1060 24618 1116
rect 24618 1060 24622 1116
rect 24558 1056 24622 1060
rect 24638 1116 24702 1120
rect 24638 1060 24642 1116
rect 24642 1060 24698 1116
rect 24698 1060 24702 1116
rect 24638 1056 24702 1060
rect 24718 1116 24782 1120
rect 24718 1060 24722 1116
rect 24722 1060 24778 1116
rect 24778 1060 24782 1116
rect 24718 1056 24782 1060
rect 32320 1116 32384 1120
rect 32320 1060 32324 1116
rect 32324 1060 32380 1116
rect 32380 1060 32384 1116
rect 32320 1056 32384 1060
rect 32400 1116 32464 1120
rect 32400 1060 32404 1116
rect 32404 1060 32460 1116
rect 32460 1060 32464 1116
rect 32400 1056 32464 1060
rect 32480 1116 32544 1120
rect 32480 1060 32484 1116
rect 32484 1060 32540 1116
rect 32540 1060 32544 1116
rect 32480 1056 32544 1060
rect 32560 1116 32624 1120
rect 32560 1060 32564 1116
rect 32564 1060 32620 1116
rect 32620 1060 32624 1116
rect 32560 1056 32624 1060
<< metal4 >>
rect 1534 17917 1594 21760
rect 2270 19549 2330 21760
rect 3006 21453 3066 21760
rect 3003 21452 3069 21453
rect 3003 21388 3004 21452
rect 3068 21388 3069 21452
rect 3003 21387 3069 21388
rect 2267 19548 2333 19549
rect 2267 19484 2268 19548
rect 2332 19484 2333 19548
rect 2267 19483 2333 19484
rect 3742 17917 3802 21760
rect 4478 21453 4538 21760
rect 5214 21453 5274 21760
rect 5950 21453 6010 21760
rect 6686 21453 6746 21760
rect 4475 21452 4541 21453
rect 4475 21388 4476 21452
rect 4540 21388 4541 21452
rect 4475 21387 4541 21388
rect 5211 21452 5277 21453
rect 5211 21388 5212 21452
rect 5276 21388 5277 21452
rect 5211 21387 5277 21388
rect 5947 21452 6013 21453
rect 5947 21388 5948 21452
rect 6012 21388 6013 21452
rect 5947 21387 6013 21388
rect 6683 21452 6749 21453
rect 6683 21388 6684 21452
rect 6748 21388 6749 21452
rect 6683 21387 6749 21388
rect 4865 20160 5185 20720
rect 7422 20637 7482 21760
rect 8158 21453 8218 21760
rect 8155 21452 8221 21453
rect 8155 21388 8156 21452
rect 8220 21388 8221 21452
rect 8155 21387 8221 21388
rect 8894 20909 8954 21760
rect 9630 21453 9690 21760
rect 9627 21452 9693 21453
rect 9627 21388 9628 21452
rect 9692 21388 9693 21452
rect 9627 21387 9693 21388
rect 10366 21317 10426 21760
rect 11102 21453 11162 21760
rect 11099 21452 11165 21453
rect 11099 21388 11100 21452
rect 11164 21388 11165 21452
rect 11099 21387 11165 21388
rect 11838 21317 11898 21760
rect 10363 21316 10429 21317
rect 10363 21252 10364 21316
rect 10428 21252 10429 21316
rect 10363 21251 10429 21252
rect 11835 21316 11901 21317
rect 11835 21252 11836 21316
rect 11900 21252 11901 21316
rect 11835 21251 11901 21252
rect 12574 21181 12634 21760
rect 12571 21180 12637 21181
rect 12571 21116 12572 21180
rect 12636 21116 12637 21180
rect 12571 21115 12637 21116
rect 8891 20908 8957 20909
rect 8891 20844 8892 20908
rect 8956 20844 8957 20908
rect 8891 20843 8957 20844
rect 8786 20704 9106 20720
rect 8786 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8954 20704
rect 9018 20640 9034 20704
rect 9098 20640 9106 20704
rect 7419 20636 7485 20637
rect 7419 20572 7420 20636
rect 7484 20572 7485 20636
rect 7419 20571 7485 20572
rect 4865 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5113 20160
rect 5177 20096 5185 20160
rect 4865 19072 5185 20096
rect 4865 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5113 19072
rect 5177 19008 5185 19072
rect 4865 17984 5185 19008
rect 4865 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5113 17984
rect 5177 17920 5185 17984
rect 1531 17916 1597 17917
rect 1531 17852 1532 17916
rect 1596 17852 1597 17916
rect 1531 17851 1597 17852
rect 3739 17916 3805 17917
rect 3739 17852 3740 17916
rect 3804 17852 3805 17916
rect 3739 17851 3805 17852
rect 4865 16896 5185 17920
rect 4865 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5113 16896
rect 5177 16832 5185 16896
rect 4865 15808 5185 16832
rect 4865 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5113 15808
rect 5177 15744 5185 15808
rect 4865 14720 5185 15744
rect 4865 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5113 14720
rect 5177 14656 5185 14720
rect 4865 13632 5185 14656
rect 4865 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5113 13632
rect 5177 13568 5185 13632
rect 4865 12544 5185 13568
rect 4865 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5113 12544
rect 5177 12480 5185 12544
rect 4865 11456 5185 12480
rect 4865 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5113 11456
rect 5177 11392 5185 11456
rect 4865 10368 5185 11392
rect 4865 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5113 10368
rect 5177 10304 5185 10368
rect 4865 9280 5185 10304
rect 4865 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5113 9280
rect 5177 9216 5185 9280
rect 4865 8192 5185 9216
rect 4865 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5113 8192
rect 5177 8128 5185 8192
rect 4865 7104 5185 8128
rect 4865 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5113 7104
rect 5177 7040 5185 7104
rect 4865 6016 5185 7040
rect 4865 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5113 6016
rect 5177 5952 5185 6016
rect 4865 4928 5185 5952
rect 4865 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5113 4928
rect 5177 4864 5185 4928
rect 4865 3840 5185 4864
rect 4865 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5113 3840
rect 5177 3776 5185 3840
rect 4865 2752 5185 3776
rect 4865 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5113 2752
rect 5177 2688 5185 2752
rect 4865 1664 5185 2688
rect 4865 1600 4873 1664
rect 4937 1600 4953 1664
rect 5017 1600 5033 1664
rect 5097 1600 5113 1664
rect 5177 1600 5185 1664
rect 4865 1040 5185 1600
rect 8786 19616 9106 20640
rect 8786 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8954 19616
rect 9018 19552 9034 19616
rect 9098 19552 9106 19616
rect 8786 18528 9106 19552
rect 8786 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8954 18528
rect 9018 18464 9034 18528
rect 9098 18464 9106 18528
rect 8786 17440 9106 18464
rect 8786 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8954 17440
rect 9018 17376 9034 17440
rect 9098 17376 9106 17440
rect 8786 16352 9106 17376
rect 8786 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8954 16352
rect 9018 16288 9034 16352
rect 9098 16288 9106 16352
rect 8786 15264 9106 16288
rect 8786 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8954 15264
rect 9018 15200 9034 15264
rect 9098 15200 9106 15264
rect 8786 14176 9106 15200
rect 8786 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8954 14176
rect 9018 14112 9034 14176
rect 9098 14112 9106 14176
rect 8786 13088 9106 14112
rect 8786 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8954 13088
rect 9018 13024 9034 13088
rect 9098 13024 9106 13088
rect 8786 12000 9106 13024
rect 8786 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8954 12000
rect 9018 11936 9034 12000
rect 9098 11936 9106 12000
rect 8786 10912 9106 11936
rect 8786 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8954 10912
rect 9018 10848 9034 10912
rect 9098 10848 9106 10912
rect 8786 9824 9106 10848
rect 8786 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8954 9824
rect 9018 9760 9034 9824
rect 9098 9760 9106 9824
rect 8786 8736 9106 9760
rect 8786 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8954 8736
rect 9018 8672 9034 8736
rect 9098 8672 9106 8736
rect 8786 7648 9106 8672
rect 8786 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8954 7648
rect 9018 7584 9034 7648
rect 9098 7584 9106 7648
rect 8786 6560 9106 7584
rect 8786 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8954 6560
rect 9018 6496 9034 6560
rect 9098 6496 9106 6560
rect 8786 5472 9106 6496
rect 8786 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8954 5472
rect 9018 5408 9034 5472
rect 9098 5408 9106 5472
rect 8786 4384 9106 5408
rect 8786 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8954 4384
rect 9018 4320 9034 4384
rect 9098 4320 9106 4384
rect 8786 3296 9106 4320
rect 8786 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8954 3296
rect 9018 3232 9034 3296
rect 9098 3232 9106 3296
rect 8786 2208 9106 3232
rect 8786 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8954 2208
rect 9018 2144 9034 2208
rect 9098 2144 9106 2208
rect 8786 1120 9106 2144
rect 8786 1056 8794 1120
rect 8858 1056 8874 1120
rect 8938 1056 8954 1120
rect 9018 1056 9034 1120
rect 9098 1056 9106 1120
rect 8786 1040 9106 1056
rect 12707 20160 13027 20720
rect 13310 20637 13370 21760
rect 14046 21453 14106 21760
rect 14782 21453 14842 21760
rect 14043 21452 14109 21453
rect 14043 21388 14044 21452
rect 14108 21388 14109 21452
rect 14043 21387 14109 21388
rect 14779 21452 14845 21453
rect 14779 21388 14780 21452
rect 14844 21388 14845 21452
rect 14779 21387 14845 21388
rect 15518 20637 15578 21760
rect 16254 21453 16314 21760
rect 16251 21452 16317 21453
rect 16251 21388 16252 21452
rect 16316 21388 16317 21452
rect 16251 21387 16317 21388
rect 16990 20909 17050 21760
rect 16987 20908 17053 20909
rect 16987 20844 16988 20908
rect 17052 20844 17053 20908
rect 16987 20843 17053 20844
rect 16628 20704 16948 20720
rect 16628 20640 16636 20704
rect 16700 20640 16716 20704
rect 16780 20640 16796 20704
rect 16860 20640 16876 20704
rect 16940 20640 16948 20704
rect 13307 20636 13373 20637
rect 13307 20572 13308 20636
rect 13372 20572 13373 20636
rect 13307 20571 13373 20572
rect 15515 20636 15581 20637
rect 15515 20572 15516 20636
rect 15580 20572 15581 20636
rect 15515 20571 15581 20572
rect 12707 20096 12715 20160
rect 12779 20096 12795 20160
rect 12859 20096 12875 20160
rect 12939 20096 12955 20160
rect 13019 20096 13027 20160
rect 12707 19072 13027 20096
rect 16628 19616 16948 20640
rect 17726 20637 17786 21760
rect 17723 20636 17789 20637
rect 17723 20572 17724 20636
rect 17788 20572 17789 20636
rect 17723 20571 17789 20572
rect 16628 19552 16636 19616
rect 16700 19552 16716 19616
rect 16780 19552 16796 19616
rect 16860 19552 16876 19616
rect 16940 19552 16948 19616
rect 13675 19412 13741 19413
rect 13675 19348 13676 19412
rect 13740 19348 13741 19412
rect 13675 19347 13741 19348
rect 12707 19008 12715 19072
rect 12779 19008 12795 19072
rect 12859 19008 12875 19072
rect 12939 19008 12955 19072
rect 13019 19008 13027 19072
rect 12707 17984 13027 19008
rect 12707 17920 12715 17984
rect 12779 17920 12795 17984
rect 12859 17920 12875 17984
rect 12939 17920 12955 17984
rect 13019 17920 13027 17984
rect 12707 16896 13027 17920
rect 12707 16832 12715 16896
rect 12779 16832 12795 16896
rect 12859 16832 12875 16896
rect 12939 16832 12955 16896
rect 13019 16832 13027 16896
rect 12707 15808 13027 16832
rect 12707 15744 12715 15808
rect 12779 15744 12795 15808
rect 12859 15744 12875 15808
rect 12939 15744 12955 15808
rect 13019 15744 13027 15808
rect 12707 14720 13027 15744
rect 12707 14656 12715 14720
rect 12779 14656 12795 14720
rect 12859 14656 12875 14720
rect 12939 14656 12955 14720
rect 13019 14656 13027 14720
rect 12707 13632 13027 14656
rect 12707 13568 12715 13632
rect 12779 13568 12795 13632
rect 12859 13568 12875 13632
rect 12939 13568 12955 13632
rect 13019 13568 13027 13632
rect 12707 12544 13027 13568
rect 12707 12480 12715 12544
rect 12779 12480 12795 12544
rect 12859 12480 12875 12544
rect 12939 12480 12955 12544
rect 13019 12480 13027 12544
rect 12707 11456 13027 12480
rect 13678 12341 13738 19347
rect 16628 18528 16948 19552
rect 18462 19549 18522 21760
rect 19198 21560 19258 21760
rect 19934 21560 19994 21760
rect 20670 21560 20730 21760
rect 21406 21560 21466 21760
rect 22142 21560 22202 21760
rect 22878 21560 22938 21760
rect 23614 21560 23674 21760
rect 24350 21560 24410 21760
rect 25086 21560 25146 21760
rect 25822 21560 25882 21760
rect 26558 21560 26618 21760
rect 27294 21045 27354 21760
rect 28030 21453 28090 21760
rect 28766 21453 28826 21760
rect 29502 21453 29562 21760
rect 28027 21452 28093 21453
rect 28027 21388 28028 21452
rect 28092 21388 28093 21452
rect 28027 21387 28093 21388
rect 28763 21452 28829 21453
rect 28763 21388 28764 21452
rect 28828 21388 28829 21452
rect 28763 21387 28829 21388
rect 29499 21452 29565 21453
rect 29499 21388 29500 21452
rect 29564 21388 29565 21452
rect 29499 21387 29565 21388
rect 27291 21044 27357 21045
rect 27291 20980 27292 21044
rect 27356 20980 27357 21044
rect 27291 20979 27357 20980
rect 20549 20160 20869 20720
rect 20549 20096 20557 20160
rect 20621 20096 20637 20160
rect 20701 20096 20717 20160
rect 20781 20096 20797 20160
rect 20861 20096 20869 20160
rect 18459 19548 18525 19549
rect 18459 19484 18460 19548
rect 18524 19484 18525 19548
rect 18459 19483 18525 19484
rect 16628 18464 16636 18528
rect 16700 18464 16716 18528
rect 16780 18464 16796 18528
rect 16860 18464 16876 18528
rect 16940 18464 16948 18528
rect 16628 17440 16948 18464
rect 16628 17376 16636 17440
rect 16700 17376 16716 17440
rect 16780 17376 16796 17440
rect 16860 17376 16876 17440
rect 16940 17376 16948 17440
rect 16628 16352 16948 17376
rect 16628 16288 16636 16352
rect 16700 16288 16716 16352
rect 16780 16288 16796 16352
rect 16860 16288 16876 16352
rect 16940 16288 16948 16352
rect 16628 15264 16948 16288
rect 16628 15200 16636 15264
rect 16700 15200 16716 15264
rect 16780 15200 16796 15264
rect 16860 15200 16876 15264
rect 16940 15200 16948 15264
rect 16628 14176 16948 15200
rect 16628 14112 16636 14176
rect 16700 14112 16716 14176
rect 16780 14112 16796 14176
rect 16860 14112 16876 14176
rect 16940 14112 16948 14176
rect 16628 13088 16948 14112
rect 16628 13024 16636 13088
rect 16700 13024 16716 13088
rect 16780 13024 16796 13088
rect 16860 13024 16876 13088
rect 16940 13024 16948 13088
rect 13675 12340 13741 12341
rect 13675 12276 13676 12340
rect 13740 12276 13741 12340
rect 13675 12275 13741 12276
rect 12707 11392 12715 11456
rect 12779 11392 12795 11456
rect 12859 11392 12875 11456
rect 12939 11392 12955 11456
rect 13019 11392 13027 11456
rect 12707 10368 13027 11392
rect 12707 10304 12715 10368
rect 12779 10304 12795 10368
rect 12859 10304 12875 10368
rect 12939 10304 12955 10368
rect 13019 10304 13027 10368
rect 12707 9280 13027 10304
rect 12707 9216 12715 9280
rect 12779 9216 12795 9280
rect 12859 9216 12875 9280
rect 12939 9216 12955 9280
rect 13019 9216 13027 9280
rect 12707 8192 13027 9216
rect 12707 8128 12715 8192
rect 12779 8128 12795 8192
rect 12859 8128 12875 8192
rect 12939 8128 12955 8192
rect 13019 8128 13027 8192
rect 12707 7104 13027 8128
rect 12707 7040 12715 7104
rect 12779 7040 12795 7104
rect 12859 7040 12875 7104
rect 12939 7040 12955 7104
rect 13019 7040 13027 7104
rect 12707 6016 13027 7040
rect 12707 5952 12715 6016
rect 12779 5952 12795 6016
rect 12859 5952 12875 6016
rect 12939 5952 12955 6016
rect 13019 5952 13027 6016
rect 12707 4928 13027 5952
rect 12707 4864 12715 4928
rect 12779 4864 12795 4928
rect 12859 4864 12875 4928
rect 12939 4864 12955 4928
rect 13019 4864 13027 4928
rect 12707 3840 13027 4864
rect 12707 3776 12715 3840
rect 12779 3776 12795 3840
rect 12859 3776 12875 3840
rect 12939 3776 12955 3840
rect 13019 3776 13027 3840
rect 12707 2752 13027 3776
rect 12707 2688 12715 2752
rect 12779 2688 12795 2752
rect 12859 2688 12875 2752
rect 12939 2688 12955 2752
rect 13019 2688 13027 2752
rect 12707 1664 13027 2688
rect 12707 1600 12715 1664
rect 12779 1600 12795 1664
rect 12859 1600 12875 1664
rect 12939 1600 12955 1664
rect 13019 1600 13027 1664
rect 12707 1040 13027 1600
rect 16628 12000 16948 13024
rect 16628 11936 16636 12000
rect 16700 11936 16716 12000
rect 16780 11936 16796 12000
rect 16860 11936 16876 12000
rect 16940 11936 16948 12000
rect 16628 10912 16948 11936
rect 16628 10848 16636 10912
rect 16700 10848 16716 10912
rect 16780 10848 16796 10912
rect 16860 10848 16876 10912
rect 16940 10848 16948 10912
rect 16628 9824 16948 10848
rect 16628 9760 16636 9824
rect 16700 9760 16716 9824
rect 16780 9760 16796 9824
rect 16860 9760 16876 9824
rect 16940 9760 16948 9824
rect 16628 8736 16948 9760
rect 16628 8672 16636 8736
rect 16700 8672 16716 8736
rect 16780 8672 16796 8736
rect 16860 8672 16876 8736
rect 16940 8672 16948 8736
rect 16628 7648 16948 8672
rect 16628 7584 16636 7648
rect 16700 7584 16716 7648
rect 16780 7584 16796 7648
rect 16860 7584 16876 7648
rect 16940 7584 16948 7648
rect 16628 6560 16948 7584
rect 16628 6496 16636 6560
rect 16700 6496 16716 6560
rect 16780 6496 16796 6560
rect 16860 6496 16876 6560
rect 16940 6496 16948 6560
rect 16628 5472 16948 6496
rect 16628 5408 16636 5472
rect 16700 5408 16716 5472
rect 16780 5408 16796 5472
rect 16860 5408 16876 5472
rect 16940 5408 16948 5472
rect 16628 4384 16948 5408
rect 16628 4320 16636 4384
rect 16700 4320 16716 4384
rect 16780 4320 16796 4384
rect 16860 4320 16876 4384
rect 16940 4320 16948 4384
rect 16628 3296 16948 4320
rect 16628 3232 16636 3296
rect 16700 3232 16716 3296
rect 16780 3232 16796 3296
rect 16860 3232 16876 3296
rect 16940 3232 16948 3296
rect 16628 2208 16948 3232
rect 16628 2144 16636 2208
rect 16700 2144 16716 2208
rect 16780 2144 16796 2208
rect 16860 2144 16876 2208
rect 16940 2144 16948 2208
rect 16628 1120 16948 2144
rect 16628 1056 16636 1120
rect 16700 1056 16716 1120
rect 16780 1056 16796 1120
rect 16860 1056 16876 1120
rect 16940 1056 16948 1120
rect 16628 1040 16948 1056
rect 20549 19072 20869 20096
rect 20549 19008 20557 19072
rect 20621 19008 20637 19072
rect 20701 19008 20717 19072
rect 20781 19008 20797 19072
rect 20861 19008 20869 19072
rect 20549 17984 20869 19008
rect 20549 17920 20557 17984
rect 20621 17920 20637 17984
rect 20701 17920 20717 17984
rect 20781 17920 20797 17984
rect 20861 17920 20869 17984
rect 20549 16896 20869 17920
rect 20549 16832 20557 16896
rect 20621 16832 20637 16896
rect 20701 16832 20717 16896
rect 20781 16832 20797 16896
rect 20861 16832 20869 16896
rect 20549 15808 20869 16832
rect 20549 15744 20557 15808
rect 20621 15744 20637 15808
rect 20701 15744 20717 15808
rect 20781 15744 20797 15808
rect 20861 15744 20869 15808
rect 20549 14720 20869 15744
rect 20549 14656 20557 14720
rect 20621 14656 20637 14720
rect 20701 14656 20717 14720
rect 20781 14656 20797 14720
rect 20861 14656 20869 14720
rect 20549 13632 20869 14656
rect 20549 13568 20557 13632
rect 20621 13568 20637 13632
rect 20701 13568 20717 13632
rect 20781 13568 20797 13632
rect 20861 13568 20869 13632
rect 20549 12544 20869 13568
rect 20549 12480 20557 12544
rect 20621 12480 20637 12544
rect 20701 12480 20717 12544
rect 20781 12480 20797 12544
rect 20861 12480 20869 12544
rect 20549 11456 20869 12480
rect 20549 11392 20557 11456
rect 20621 11392 20637 11456
rect 20701 11392 20717 11456
rect 20781 11392 20797 11456
rect 20861 11392 20869 11456
rect 20549 10368 20869 11392
rect 20549 10304 20557 10368
rect 20621 10304 20637 10368
rect 20701 10304 20717 10368
rect 20781 10304 20797 10368
rect 20861 10304 20869 10368
rect 20549 9280 20869 10304
rect 20549 9216 20557 9280
rect 20621 9216 20637 9280
rect 20701 9216 20717 9280
rect 20781 9216 20797 9280
rect 20861 9216 20869 9280
rect 20549 8192 20869 9216
rect 20549 8128 20557 8192
rect 20621 8128 20637 8192
rect 20701 8128 20717 8192
rect 20781 8128 20797 8192
rect 20861 8128 20869 8192
rect 20549 7104 20869 8128
rect 20549 7040 20557 7104
rect 20621 7040 20637 7104
rect 20701 7040 20717 7104
rect 20781 7040 20797 7104
rect 20861 7040 20869 7104
rect 20549 6016 20869 7040
rect 20549 5952 20557 6016
rect 20621 5952 20637 6016
rect 20701 5952 20717 6016
rect 20781 5952 20797 6016
rect 20861 5952 20869 6016
rect 20549 4928 20869 5952
rect 20549 4864 20557 4928
rect 20621 4864 20637 4928
rect 20701 4864 20717 4928
rect 20781 4864 20797 4928
rect 20861 4864 20869 4928
rect 20549 3840 20869 4864
rect 20549 3776 20557 3840
rect 20621 3776 20637 3840
rect 20701 3776 20717 3840
rect 20781 3776 20797 3840
rect 20861 3776 20869 3840
rect 20549 2752 20869 3776
rect 20549 2688 20557 2752
rect 20621 2688 20637 2752
rect 20701 2688 20717 2752
rect 20781 2688 20797 2752
rect 20861 2688 20869 2752
rect 20549 1664 20869 2688
rect 20549 1600 20557 1664
rect 20621 1600 20637 1664
rect 20701 1600 20717 1664
rect 20781 1600 20797 1664
rect 20861 1600 20869 1664
rect 20549 1040 20869 1600
rect 24470 20704 24790 20720
rect 24470 20640 24478 20704
rect 24542 20640 24558 20704
rect 24622 20640 24638 20704
rect 24702 20640 24718 20704
rect 24782 20640 24790 20704
rect 24470 19616 24790 20640
rect 24470 19552 24478 19616
rect 24542 19552 24558 19616
rect 24622 19552 24638 19616
rect 24702 19552 24718 19616
rect 24782 19552 24790 19616
rect 24470 18528 24790 19552
rect 24470 18464 24478 18528
rect 24542 18464 24558 18528
rect 24622 18464 24638 18528
rect 24702 18464 24718 18528
rect 24782 18464 24790 18528
rect 24470 17440 24790 18464
rect 24470 17376 24478 17440
rect 24542 17376 24558 17440
rect 24622 17376 24638 17440
rect 24702 17376 24718 17440
rect 24782 17376 24790 17440
rect 24470 16352 24790 17376
rect 24470 16288 24478 16352
rect 24542 16288 24558 16352
rect 24622 16288 24638 16352
rect 24702 16288 24718 16352
rect 24782 16288 24790 16352
rect 24470 15264 24790 16288
rect 24470 15200 24478 15264
rect 24542 15200 24558 15264
rect 24622 15200 24638 15264
rect 24702 15200 24718 15264
rect 24782 15200 24790 15264
rect 24470 14176 24790 15200
rect 24470 14112 24478 14176
rect 24542 14112 24558 14176
rect 24622 14112 24638 14176
rect 24702 14112 24718 14176
rect 24782 14112 24790 14176
rect 24470 13088 24790 14112
rect 24470 13024 24478 13088
rect 24542 13024 24558 13088
rect 24622 13024 24638 13088
rect 24702 13024 24718 13088
rect 24782 13024 24790 13088
rect 24470 12000 24790 13024
rect 24470 11936 24478 12000
rect 24542 11936 24558 12000
rect 24622 11936 24638 12000
rect 24702 11936 24718 12000
rect 24782 11936 24790 12000
rect 24470 10912 24790 11936
rect 24470 10848 24478 10912
rect 24542 10848 24558 10912
rect 24622 10848 24638 10912
rect 24702 10848 24718 10912
rect 24782 10848 24790 10912
rect 24470 9824 24790 10848
rect 24470 9760 24478 9824
rect 24542 9760 24558 9824
rect 24622 9760 24638 9824
rect 24702 9760 24718 9824
rect 24782 9760 24790 9824
rect 24470 8736 24790 9760
rect 24470 8672 24478 8736
rect 24542 8672 24558 8736
rect 24622 8672 24638 8736
rect 24702 8672 24718 8736
rect 24782 8672 24790 8736
rect 24470 7648 24790 8672
rect 24470 7584 24478 7648
rect 24542 7584 24558 7648
rect 24622 7584 24638 7648
rect 24702 7584 24718 7648
rect 24782 7584 24790 7648
rect 24470 6560 24790 7584
rect 24470 6496 24478 6560
rect 24542 6496 24558 6560
rect 24622 6496 24638 6560
rect 24702 6496 24718 6560
rect 24782 6496 24790 6560
rect 24470 5472 24790 6496
rect 24470 5408 24478 5472
rect 24542 5408 24558 5472
rect 24622 5408 24638 5472
rect 24702 5408 24718 5472
rect 24782 5408 24790 5472
rect 24470 4384 24790 5408
rect 24470 4320 24478 4384
rect 24542 4320 24558 4384
rect 24622 4320 24638 4384
rect 24702 4320 24718 4384
rect 24782 4320 24790 4384
rect 24470 3296 24790 4320
rect 24470 3232 24478 3296
rect 24542 3232 24558 3296
rect 24622 3232 24638 3296
rect 24702 3232 24718 3296
rect 24782 3232 24790 3296
rect 24470 2208 24790 3232
rect 24470 2144 24478 2208
rect 24542 2144 24558 2208
rect 24622 2144 24638 2208
rect 24702 2144 24718 2208
rect 24782 2144 24790 2208
rect 24470 1120 24790 2144
rect 24470 1056 24478 1120
rect 24542 1056 24558 1120
rect 24622 1056 24638 1120
rect 24702 1056 24718 1120
rect 24782 1056 24790 1120
rect 24470 1040 24790 1056
rect 28391 20160 28711 20720
rect 28391 20096 28399 20160
rect 28463 20096 28479 20160
rect 28543 20096 28559 20160
rect 28623 20096 28639 20160
rect 28703 20096 28711 20160
rect 28391 19072 28711 20096
rect 28391 19008 28399 19072
rect 28463 19008 28479 19072
rect 28543 19008 28559 19072
rect 28623 19008 28639 19072
rect 28703 19008 28711 19072
rect 28391 17984 28711 19008
rect 28391 17920 28399 17984
rect 28463 17920 28479 17984
rect 28543 17920 28559 17984
rect 28623 17920 28639 17984
rect 28703 17920 28711 17984
rect 28391 16896 28711 17920
rect 30238 16965 30298 21760
rect 30974 21453 31034 21760
rect 30971 21452 31037 21453
rect 30971 21388 30972 21452
rect 31036 21388 31037 21452
rect 31710 21450 31770 21760
rect 32446 21560 32506 21760
rect 30971 21387 31037 21388
rect 31526 21390 31770 21450
rect 31526 17917 31586 21390
rect 32312 20704 32632 20720
rect 32312 20640 32320 20704
rect 32384 20640 32400 20704
rect 32464 20640 32480 20704
rect 32544 20640 32560 20704
rect 32624 20640 32632 20704
rect 32312 19616 32632 20640
rect 32312 19552 32320 19616
rect 32384 19552 32400 19616
rect 32464 19552 32480 19616
rect 32544 19552 32560 19616
rect 32624 19552 32632 19616
rect 32312 18528 32632 19552
rect 32312 18464 32320 18528
rect 32384 18464 32400 18528
rect 32464 18464 32480 18528
rect 32544 18464 32560 18528
rect 32624 18464 32632 18528
rect 31523 17916 31589 17917
rect 31523 17852 31524 17916
rect 31588 17852 31589 17916
rect 31523 17851 31589 17852
rect 32312 17440 32632 18464
rect 32312 17376 32320 17440
rect 32384 17376 32400 17440
rect 32464 17376 32480 17440
rect 32544 17376 32560 17440
rect 32624 17376 32632 17440
rect 30235 16964 30301 16965
rect 30235 16900 30236 16964
rect 30300 16900 30301 16964
rect 30235 16899 30301 16900
rect 28391 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28639 16896
rect 28703 16832 28711 16896
rect 28391 15808 28711 16832
rect 28391 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28639 15808
rect 28703 15744 28711 15808
rect 28391 14720 28711 15744
rect 28391 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28639 14720
rect 28703 14656 28711 14720
rect 28391 13632 28711 14656
rect 28391 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28639 13632
rect 28703 13568 28711 13632
rect 28391 12544 28711 13568
rect 28391 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28639 12544
rect 28703 12480 28711 12544
rect 28391 11456 28711 12480
rect 28391 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28639 11456
rect 28703 11392 28711 11456
rect 28391 10368 28711 11392
rect 28391 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28639 10368
rect 28703 10304 28711 10368
rect 28391 9280 28711 10304
rect 28391 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28639 9280
rect 28703 9216 28711 9280
rect 28391 8192 28711 9216
rect 28391 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28639 8192
rect 28703 8128 28711 8192
rect 28391 7104 28711 8128
rect 28391 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28639 7104
rect 28703 7040 28711 7104
rect 28391 6016 28711 7040
rect 28391 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28639 6016
rect 28703 5952 28711 6016
rect 28391 4928 28711 5952
rect 28391 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28639 4928
rect 28703 4864 28711 4928
rect 28391 3840 28711 4864
rect 28391 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28639 3840
rect 28703 3776 28711 3840
rect 28391 2752 28711 3776
rect 28391 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28639 2752
rect 28703 2688 28711 2752
rect 28391 1664 28711 2688
rect 28391 1600 28399 1664
rect 28463 1600 28479 1664
rect 28543 1600 28559 1664
rect 28623 1600 28639 1664
rect 28703 1600 28711 1664
rect 28391 1040 28711 1600
rect 32312 16352 32632 17376
rect 32312 16288 32320 16352
rect 32384 16288 32400 16352
rect 32464 16288 32480 16352
rect 32544 16288 32560 16352
rect 32624 16288 32632 16352
rect 32312 15264 32632 16288
rect 32312 15200 32320 15264
rect 32384 15200 32400 15264
rect 32464 15200 32480 15264
rect 32544 15200 32560 15264
rect 32624 15200 32632 15264
rect 32312 14176 32632 15200
rect 32312 14112 32320 14176
rect 32384 14112 32400 14176
rect 32464 14112 32480 14176
rect 32544 14112 32560 14176
rect 32624 14112 32632 14176
rect 32312 13088 32632 14112
rect 32312 13024 32320 13088
rect 32384 13024 32400 13088
rect 32464 13024 32480 13088
rect 32544 13024 32560 13088
rect 32624 13024 32632 13088
rect 32312 12000 32632 13024
rect 32312 11936 32320 12000
rect 32384 11936 32400 12000
rect 32464 11936 32480 12000
rect 32544 11936 32560 12000
rect 32624 11936 32632 12000
rect 32312 10912 32632 11936
rect 32312 10848 32320 10912
rect 32384 10848 32400 10912
rect 32464 10848 32480 10912
rect 32544 10848 32560 10912
rect 32624 10848 32632 10912
rect 32312 9824 32632 10848
rect 32312 9760 32320 9824
rect 32384 9760 32400 9824
rect 32464 9760 32480 9824
rect 32544 9760 32560 9824
rect 32624 9760 32632 9824
rect 32312 8736 32632 9760
rect 32312 8672 32320 8736
rect 32384 8672 32400 8736
rect 32464 8672 32480 8736
rect 32544 8672 32560 8736
rect 32624 8672 32632 8736
rect 32312 7648 32632 8672
rect 32312 7584 32320 7648
rect 32384 7584 32400 7648
rect 32464 7584 32480 7648
rect 32544 7584 32560 7648
rect 32624 7584 32632 7648
rect 32312 6560 32632 7584
rect 32312 6496 32320 6560
rect 32384 6496 32400 6560
rect 32464 6496 32480 6560
rect 32544 6496 32560 6560
rect 32624 6496 32632 6560
rect 32312 5472 32632 6496
rect 32312 5408 32320 5472
rect 32384 5408 32400 5472
rect 32464 5408 32480 5472
rect 32544 5408 32560 5472
rect 32624 5408 32632 5472
rect 32312 4384 32632 5408
rect 32312 4320 32320 4384
rect 32384 4320 32400 4384
rect 32464 4320 32480 4384
rect 32544 4320 32560 4384
rect 32624 4320 32632 4384
rect 32312 3296 32632 4320
rect 32312 3232 32320 3296
rect 32384 3232 32400 3296
rect 32464 3232 32480 3296
rect 32544 3232 32560 3296
rect 32624 3232 32632 3296
rect 32312 2208 32632 3232
rect 32312 2144 32320 2208
rect 32384 2144 32400 2208
rect 32464 2144 32480 2208
rect 32544 2144 32560 2208
rect 32624 2144 32632 2208
rect 32312 1120 32632 2144
rect 32312 1056 32320 1120
rect 32384 1056 32400 1120
rect 32464 1056 32480 1120
rect 32544 1056 32560 1120
rect 32624 1056 32632 1120
rect 32312 1040 32632 1056
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_337
timestamp 1676037725
transform 1 0 32108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_337
timestamp 1676037725
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_174
timestamp 1676037725
transform 1 0 17112 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_198 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_206
timestamp 1676037725
transform 1 0 20056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_213
timestamp 1676037725
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1676037725
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_127
timestamp 1676037725
transform 1 0 12788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_161
timestamp 1676037725
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1676037725
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1676037725
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1676037725
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_205
timestamp 1676037725
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_214
timestamp 1676037725
transform 1 0 20792 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_224
timestamp 1676037725
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_234
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1676037725
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_337
timestamp 1676037725
transform 1 0 32108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1676037725
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1676037725
transform 1 0 8096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_92
timestamp 1676037725
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1676037725
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_117
timestamp 1676037725
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1676037725
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_135
timestamp 1676037725
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_147
timestamp 1676037725
transform 1 0 14628 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1676037725
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1676037725
transform 1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1676037725
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1676037725
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_233
timestamp 1676037725
transform 1 0 22540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_245
timestamp 1676037725
transform 1 0 23644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_257
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1676037725
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1676037725
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_35
timestamp 1676037725
transform 1 0 4324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1676037725
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1676037725
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_58
timestamp 1676037725
transform 1 0 6440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_62
timestamp 1676037725
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1676037725
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp 1676037725
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_102
timestamp 1676037725
transform 1 0 10488 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1676037725
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1676037725
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_149
timestamp 1676037725
transform 1 0 14812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1676037725
transform 1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_203
timestamp 1676037725
transform 1 0 19780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_217
timestamp 1676037725
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_227
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_242
timestamp 1676037725
transform 1 0 23368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1676037725
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_337
timestamp 1676037725
transform 1 0 32108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1676037725
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_45
timestamp 1676037725
transform 1 0 5244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1676037725
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_72
timestamp 1676037725
transform 1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_82
timestamp 1676037725
transform 1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1676037725
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1676037725
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_128
timestamp 1676037725
transform 1 0 12880 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_150
timestamp 1676037725
transform 1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_183
timestamp 1676037725
transform 1 0 17940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_195
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1676037725
transform 1 0 19780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_210
timestamp 1676037725
transform 1 0 20424 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1676037725
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_236
timestamp 1676037725
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1676037725
transform 1 0 24840 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_266
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1676037725
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1676037725
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1676037725
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_100
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_108
timestamp 1676037725
transform 1 0 11040 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_112
timestamp 1676037725
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1676037725
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1676037725
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_180
timestamp 1676037725
transform 1 0 17664 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1676037725
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_214
timestamp 1676037725
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_239
timestamp 1676037725
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1676037725
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_282
timestamp 1676037725
transform 1 0 27048 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_293
timestamp 1676037725
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1676037725
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_337
timestamp 1676037725
transform 1 0 32108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1676037725
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1676037725
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1676037725
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_63
timestamp 1676037725
transform 1 0 6900 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_84
timestamp 1676037725
transform 1 0 8832 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1676037725
transform 1 0 9568 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1676037725
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1676037725
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1676037725
transform 1 0 12420 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 1676037725
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_131
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_144
timestamp 1676037725
transform 1 0 14352 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_192
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_247
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_254
timestamp 1676037725
transform 1 0 24472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_260
timestamp 1676037725
transform 1 0 25024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_300
timestamp 1676037725
transform 1 0 28704 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_308
timestamp 1676037725
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_326
timestamp 1676037725
transform 1 0 31096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1676037725
transform 1 0 4416 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_52
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1676037725
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_75
timestamp 1676037725
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_98
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_120
timestamp 1676037725
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_168
timestamp 1676037725
transform 1 0 16560 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_180
timestamp 1676037725
transform 1 0 17664 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_188
timestamp 1676037725
transform 1 0 18400 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1676037725
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_223
timestamp 1676037725
transform 1 0 21620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_260
timestamp 1676037725
transform 1 0 25024 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_273
timestamp 1676037725
transform 1 0 26220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1676037725
transform 1 0 27232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_297
timestamp 1676037725
transform 1 0 28428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1676037725
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_337
timestamp 1676037725
transform 1 0 32108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1676037725
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1676037725
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_40
timestamp 1676037725
transform 1 0 4784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_48
timestamp 1676037725
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_80
timestamp 1676037725
transform 1 0 8464 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_88
timestamp 1676037725
transform 1 0 9200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1676037725
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_155
timestamp 1676037725
transform 1 0 15364 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_191
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_250
timestamp 1676037725
transform 1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_258
timestamp 1676037725
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1676037725
transform 1 0 25760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_272
timestamp 1676037725
transform 1 0 26128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1676037725
transform 1 0 28980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_311
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1676037725
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1676037725
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1676037725
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1676037725
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1676037725
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1676037725
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1676037725
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1676037725
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_158
timestamp 1676037725
transform 1 0 15640 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1676037725
transform 1 0 16192 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_234
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_243
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 1676037725
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_266
timestamp 1676037725
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_290
timestamp 1676037725
transform 1 0 27784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_319
timestamp 1676037725
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_329
timestamp 1676037725
transform 1 0 31372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_336
timestamp 1676037725
transform 1 0 32016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_28
timestamp 1676037725
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1676037725
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_118
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_126
timestamp 1676037725
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_178
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1676037725
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1676037725
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_235
timestamp 1676037725
transform 1 0 22724 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_241
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1676037725
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1676037725
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1676037725
transform 1 0 29256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1676037725
transform 1 0 30084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_323
timestamp 1676037725
transform 1 0 30820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1676037725
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_35
timestamp 1676037725
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1676037725
transform 1 0 5152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1676037725
transform 1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1676037725
transform 1 0 8280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_100
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_104
timestamp 1676037725
transform 1 0 10672 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_116
timestamp 1676037725
transform 1 0 11776 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_160
timestamp 1676037725
transform 1 0 15824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_220
timestamp 1676037725
transform 1 0 21344 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_232
timestamp 1676037725
transform 1 0 22448 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1676037725
transform 1 0 23184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_262
timestamp 1676037725
transform 1 0 25208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_266
timestamp 1676037725
transform 1 0 25576 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1676037725
transform 1 0 26128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_280
timestamp 1676037725
transform 1 0 26864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_295
timestamp 1676037725
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_299
timestamp 1676037725
transform 1 0 28612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_317
timestamp 1676037725
transform 1 0 30268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_329
timestamp 1676037725
transform 1 0 31372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_337
timestamp 1676037725
transform 1 0 32108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1676037725
transform 1 0 3496 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_65
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_77
timestamp 1676037725
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_133
timestamp 1676037725
transform 1 0 13340 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_160
timestamp 1676037725
transform 1 0 15824 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_186
timestamp 1676037725
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_196
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1676037725
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_234
timestamp 1676037725
transform 1 0 22632 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1676037725
transform 1 0 23368 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_247
timestamp 1676037725
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_259
timestamp 1676037725
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_271
timestamp 1676037725
transform 1 0 26036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1676037725
transform 1 0 27508 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_299
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_308
timestamp 1676037725
transform 1 0 29440 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_315
timestamp 1676037725
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_326
timestamp 1676037725
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_35
timestamp 1676037725
transform 1 0 4324 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_47
timestamp 1676037725
transform 1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1676037725
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_67
timestamp 1676037725
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1676037725
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1676037725
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_171
timestamp 1676037725
transform 1 0 16836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_223
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1676037725
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_243
timestamp 1676037725
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1676037725
transform 1 0 25208 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_275
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_287
timestamp 1676037725
transform 1 0 27508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_298
timestamp 1676037725
transform 1 0 28520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1676037725
transform 1 0 30360 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_325
timestamp 1676037725
transform 1 0 31004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_337
timestamp 1676037725
transform 1 0 32108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_36
timestamp 1676037725
transform 1 0 4416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_43
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_77
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_94
timestamp 1676037725
transform 1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1676037725
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_215
timestamp 1676037725
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_236
timestamp 1676037725
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_248
timestamp 1676037725
transform 1 0 23920 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_257
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_265
timestamp 1676037725
transform 1 0 25484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_289
timestamp 1676037725
transform 1 0 27692 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_300
timestamp 1676037725
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_313
timestamp 1676037725
transform 1 0 29900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1676037725
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1676037725
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_36
timestamp 1676037725
transform 1 0 4416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1676037725
transform 1 0 4784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1676037725
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1676037725
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_114
timestamp 1676037725
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_127
timestamp 1676037725
transform 1 0 12788 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1676037725
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_157
timestamp 1676037725
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_169
timestamp 1676037725
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_203
timestamp 1676037725
transform 1 0 19780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_258
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_274
timestamp 1676037725
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1676037725
transform 1 0 26956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1676037725
transform 1 0 28520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_318
timestamp 1676037725
transform 1 0 30360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_330
timestamp 1676037725
transform 1 0 31464 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1676037725
transform 1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_31
timestamp 1676037725
transform 1 0 3956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_42
timestamp 1676037725
transform 1 0 4968 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1676037725
transform 1 0 5520 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1676037725
transform 1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_79
timestamp 1676037725
transform 1 0 8372 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1676037725
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_118
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_130
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1676037725
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1676037725
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1676037725
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_242
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_250
timestamp 1676037725
transform 1 0 24104 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_255
timestamp 1676037725
transform 1 0 24564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_270
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1676037725
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1676037725
transform 1 0 29900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_322
timestamp 1676037725
transform 1 0 30728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_36
timestamp 1676037725
transform 1 0 4416 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_48
timestamp 1676037725
transform 1 0 5520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1676037725
transform 1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1676037725
transform 1 0 6808 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1676037725
transform 1 0 8004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1676037725
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1676037725
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_274
timestamp 1676037725
transform 1 0 26312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_282
timestamp 1676037725
transform 1 0 27048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_290
timestamp 1676037725
transform 1 0 27784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_296
timestamp 1676037725
transform 1 0 28336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1676037725
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_328
timestamp 1676037725
transform 1 0 31280 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_336
timestamp 1676037725
transform 1 0 32016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1676037725
transform 1 0 2944 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_31
timestamp 1676037725
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_43
timestamp 1676037725
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_67
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1676037725
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1676037725
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1676037725
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1676037725
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_241
timestamp 1676037725
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_288
timestamp 1676037725
transform 1 0 27600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_297
timestamp 1676037725
transform 1 0 28428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_313
timestamp 1676037725
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1676037725
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_8
timestamp 1676037725
transform 1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_19
timestamp 1676037725
transform 1 0 2852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1676037725
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1676037725
transform 1 0 11960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_127
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_184
timestamp 1676037725
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_188
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1676037725
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_212
timestamp 1676037725
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1676037725
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_259
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_267
timestamp 1676037725
transform 1 0 25668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1676037725
transform 1 0 27876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_302
timestamp 1676037725
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_314
timestamp 1676037725
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_328
timestamp 1676037725
transform 1 0 31280 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_336
timestamp 1676037725
transform 1 0 32016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_8
timestamp 1676037725
transform 1 0 1840 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_14
timestamp 1676037725
transform 1 0 2392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_22
timestamp 1676037725
transform 1 0 3128 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_30
timestamp 1676037725
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_37
timestamp 1676037725
transform 1 0 4508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_41
timestamp 1676037725
transform 1 0 4876 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_46
timestamp 1676037725
transform 1 0 5336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_65
timestamp 1676037725
transform 1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp 1676037725
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_121
timestamp 1676037725
transform 1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_177
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1676037725
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1676037725
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_257
timestamp 1676037725
transform 1 0 24748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1676037725
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_294
timestamp 1676037725
transform 1 0 28152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_299
timestamp 1676037725
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1676037725
transform 1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_327
timestamp 1676037725
transform 1 0 31188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_14
timestamp 1676037725
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1676037725
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_48
timestamp 1676037725
transform 1 0 5520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_76
timestamp 1676037725
transform 1 0 8096 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1676037725
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_107
timestamp 1676037725
transform 1 0 10948 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_115
timestamp 1676037725
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_120
timestamp 1676037725
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1676037725
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1676037725
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1676037725
transform 1 0 16008 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1676037725
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_261
timestamp 1676037725
transform 1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_269
timestamp 1676037725
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_291
timestamp 1676037725
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_327
timestamp 1676037725
transform 1 0 31188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_335
timestamp 1676037725
transform 1 0 31924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_16
timestamp 1676037725
transform 1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_25
timestamp 1676037725
transform 1 0 3404 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1676037725
transform 1 0 3956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_48
timestamp 1676037725
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1676037725
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_67
timestamp 1676037725
transform 1 0 7268 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_102
timestamp 1676037725
transform 1 0 10488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1676037725
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1676037725
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_140
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_155
timestamp 1676037725
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_177
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_183
timestamp 1676037725
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 1676037725
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_230
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_238
timestamp 1676037725
transform 1 0 23000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_255
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_266
timestamp 1676037725
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_270
timestamp 1676037725
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_285
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_302
timestamp 1676037725
transform 1 0 28888 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_308
timestamp 1676037725
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1676037725
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1676037725
transform 1 0 2576 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1676037725
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_49
timestamp 1676037725
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_66
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1676037725
transform 1 0 11776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_128
timestamp 1676037725
transform 1 0 12880 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_132
timestamp 1676037725
transform 1 0 13248 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_155
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_168
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_174
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_182
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_206
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_218
timestamp 1676037725
transform 1 0 21160 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_230
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_261
timestamp 1676037725
transform 1 0 25116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_267
timestamp 1676037725
transform 1 0 25668 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1676037725
transform 1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_329
timestamp 1676037725
transform 1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_336
timestamp 1676037725
transform 1 0 32016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1676037725
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_17
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_63
timestamp 1676037725
transform 1 0 6900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_80
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_88
timestamp 1676037725
transform 1 0 9200 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_94
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1676037725
transform 1 0 10212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 1676037725
transform 1 0 10580 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_127
timestamp 1676037725
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_203
timestamp 1676037725
transform 1 0 19780 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_213
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_230
timestamp 1676037725
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_245
timestamp 1676037725
transform 1 0 23644 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1676037725
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_257
timestamp 1676037725
transform 1 0 24748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_287
timestamp 1676037725
transform 1 0 27508 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_291
timestamp 1676037725
transform 1 0 27876 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_300
timestamp 1676037725
transform 1 0 28704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_320
timestamp 1676037725
transform 1 0 30544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_14
timestamp 1676037725
transform 1 0 2392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1676037725
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_39
timestamp 1676037725
transform 1 0 4692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_50
timestamp 1676037725
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1676037725
transform 1 0 6348 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_95
timestamp 1676037725
transform 1 0 9844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_103
timestamp 1676037725
transform 1 0 10580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1676037725
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1676037725
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_219
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_232
timestamp 1676037725
transform 1 0 22448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1676037725
transform 1 0 23184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_269
timestamp 1676037725
transform 1 0 25852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_287
timestamp 1676037725
transform 1 0 27508 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_300
timestamp 1676037725
transform 1 0 28704 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1676037725
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_328
timestamp 1676037725
transform 1 0 31280 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_335
timestamp 1676037725
transform 1 0 31924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_8
timestamp 1676037725
transform 1 0 1840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_25
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_65
timestamp 1676037725
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1676037725
transform 1 0 7912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_83
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_100
timestamp 1676037725
transform 1 0 10304 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_139
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_175
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1676037725
transform 1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_234
timestamp 1676037725
transform 1 0 22632 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_245
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_256
timestamp 1676037725
transform 1 0 24656 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1676037725
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_290
timestamp 1676037725
transform 1 0 27784 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_312
timestamp 1676037725
transform 1 0 29808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_12
timestamp 1676037725
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_19
timestamp 1676037725
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_48
timestamp 1676037725
transform 1 0 5520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_55
timestamp 1676037725
transform 1 0 6164 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_63
timestamp 1676037725
transform 1 0 6900 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_104
timestamp 1676037725
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_111
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_132
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1676037725
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_218
timestamp 1676037725
transform 1 0 21160 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_226
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1676037725
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_266
timestamp 1676037725
transform 1 0 25576 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1676037725
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_281
timestamp 1676037725
transform 1 0 26956 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1676037725
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1676037725
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_335
timestamp 1676037725
transform 1 0 31924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_12
timestamp 1676037725
transform 1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_19
timestamp 1676037725
transform 1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_26
timestamp 1676037725
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_29
timestamp 1676037725
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_43
timestamp 1676037725
transform 1 0 5060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_62
timestamp 1676037725
transform 1 0 6808 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_71
timestamp 1676037725
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_79
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_83
timestamp 1676037725
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1676037725
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_89
timestamp 1676037725
transform 1 0 9292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_94
timestamp 1676037725
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1676037725
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1676037725
transform 1 0 13248 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_141
timestamp 1676037725
transform 1 0 14076 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_175
timestamp 1676037725
transform 1 0 17204 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_212
timestamp 1676037725
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_246
timestamp 1676037725
transform 1 0 23736 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1676037725
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_294
timestamp 1676037725
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_306
timestamp 1676037725
transform 1 0 29256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_309
timestamp 1676037725
transform 1 0 29532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_327
timestamp 1676037725
transform 1 0 31188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 32476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 32476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 32476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 32476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 32476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 32476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 32476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 32476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 32476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 32476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 32476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 32476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 32476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 32476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 32476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 32476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 32476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 32476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 32476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 32476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 32476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 32476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 32476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 32476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 32476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 32476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 32476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 32476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 32476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 32476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 32476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 32476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 32476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15364 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0503_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0505_
timestamp 1676037725
transform -1 0 25576 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0506_
timestamp 1676037725
transform 1 0 14536 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8280 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _0512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0514_
timestamp 1676037725
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0515_
timestamp 1676037725
transform 1 0 20976 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0517_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0518_
timestamp 1676037725
transform -1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0519_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1676037725
transform -1 0 14352 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _0521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11776 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0522_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12788 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0523_
timestamp 1676037725
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0524_
timestamp 1676037725
transform 1 0 10764 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0525_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11592 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0530_
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0532_
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0533_
timestamp 1676037725
transform -1 0 8280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0535_
timestamp 1676037725
transform -1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13984 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0537_
timestamp 1676037725
transform -1 0 25116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1676037725
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0539_
timestamp 1676037725
transform -1 0 27508 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0540_
timestamp 1676037725
transform -1 0 24012 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0541_
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1676037725
transform -1 0 5704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0543_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0544_
timestamp 1676037725
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0545_
timestamp 1676037725
transform 1 0 13156 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1676037725
transform -1 0 25484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0548_
timestamp 1676037725
transform 1 0 15732 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16560 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12328 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_4  _0551_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13892 0 -1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__o32a_1  _0552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12512 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0554_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12144 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0556_
timestamp 1676037725
transform -1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1676037725
transform -1 0 7636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0560_
timestamp 1676037725
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0561_
timestamp 1676037725
transform -1 0 20240 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1676037725
transform -1 0 6348 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0564_
timestamp 1676037725
transform -1 0 17848 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0565_
timestamp 1676037725
transform -1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0566_
timestamp 1676037725
transform -1 0 17940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0567_
timestamp 1676037725
transform -1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10028 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0571_
timestamp 1676037725
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0572_
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0573_
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0574_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0575_
timestamp 1676037725
transform 1 0 16376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0576_
timestamp 1676037725
transform -1 0 16008 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27508 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1676037725
transform -1 0 8648 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0579_
timestamp 1676037725
transform 1 0 24472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0580_
timestamp 1676037725
transform -1 0 20792 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0581_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0582_
timestamp 1676037725
transform -1 0 20056 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0583_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23644 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0585_
timestamp 1676037725
transform -1 0 26404 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26128 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0587_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0588_
timestamp 1676037725
transform 1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0589_
timestamp 1676037725
transform 1 0 19412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0590_
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0591_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0593_
timestamp 1676037725
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0594_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0596_
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0597_
timestamp 1676037725
transform -1 0 23276 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0598_
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0599_
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0600_
timestamp 1676037725
transform -1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0601_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0602_
timestamp 1676037725
transform 1 0 20332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0603_
timestamp 1676037725
transform 1 0 21988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0605_
timestamp 1676037725
transform -1 0 20884 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0606_
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0607_
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0608_
timestamp 1676037725
transform 1 0 25944 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0609_
timestamp 1676037725
transform 1 0 25852 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0610_
timestamp 1676037725
transform -1 0 27784 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0611_
timestamp 1676037725
transform -1 0 26956 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0612_
timestamp 1676037725
transform 1 0 24012 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0613_
timestamp 1676037725
transform -1 0 25208 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0615_
timestamp 1676037725
transform -1 0 16284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0616_
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0619_
timestamp 1676037725
transform -1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _0622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0623_
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0624_
timestamp 1676037725
transform -1 0 20332 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0625_
timestamp 1676037725
transform -1 0 17756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0626_
timestamp 1676037725
transform -1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0627_
timestamp 1676037725
transform 1 0 2944 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0628_
timestamp 1676037725
transform -1 0 3404 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0629_
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1676037725
transform -1 0 3496 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0632_
timestamp 1676037725
transform 1 0 27784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1676037725
transform 1 0 31556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0634_
timestamp 1676037725
transform -1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0635_
timestamp 1676037725
transform -1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0636_
timestamp 1676037725
transform 1 0 15088 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0637_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0638_
timestamp 1676037725
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0639_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0640_
timestamp 1676037725
transform -1 0 6992 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0641_
timestamp 1676037725
transform -1 0 15916 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14904 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0643_
timestamp 1676037725
transform -1 0 8464 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0646_
timestamp 1676037725
transform -1 0 29256 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0647_
timestamp 1676037725
transform 1 0 21712 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0648_
timestamp 1676037725
transform -1 0 25116 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0649_
timestamp 1676037725
transform -1 0 24564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0650_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1676037725
transform 1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0652_
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14720 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0654_
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0655_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1676037725
transform -1 0 31924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0657_
timestamp 1676037725
transform -1 0 25116 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22724 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0659_
timestamp 1676037725
transform -1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0660_
timestamp 1676037725
transform -1 0 8372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0661_
timestamp 1676037725
transform -1 0 7912 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0662_
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0664_
timestamp 1676037725
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0665_
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0666_
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0668_
timestamp 1676037725
transform -1 0 23920 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0669_
timestamp 1676037725
transform -1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0670_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0672_
timestamp 1676037725
transform -1 0 22540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0673_
timestamp 1676037725
transform -1 0 22632 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23920 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0675_
timestamp 1676037725
transform -1 0 21988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0676_
timestamp 1676037725
transform -1 0 21436 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0677_
timestamp 1676037725
transform -1 0 22816 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0678_
timestamp 1676037725
transform -1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0679_
timestamp 1676037725
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0680_
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1676037725
transform -1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0682_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0683_
timestamp 1676037725
transform -1 0 24196 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23736 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _0685_
timestamp 1676037725
transform 1 0 20240 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0686_
timestamp 1676037725
transform 1 0 19596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0687_
timestamp 1676037725
transform 1 0 20424 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _0688_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21160 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0689_
timestamp 1676037725
transform -1 0 20424 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0690_
timestamp 1676037725
transform -1 0 19964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0691_
timestamp 1676037725
transform -1 0 18492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0692_
timestamp 1676037725
transform -1 0 17664 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0694_
timestamp 1676037725
transform 1 0 20148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0695_
timestamp 1676037725
transform 1 0 20792 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0696_
timestamp 1676037725
transform 1 0 20516 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0697_
timestamp 1676037725
transform 1 0 16836 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0698_
timestamp 1676037725
transform -1 0 17940 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0699_
timestamp 1676037725
transform -1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0700_
timestamp 1676037725
transform 1 0 14720 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0701_
timestamp 1676037725
transform 1 0 15916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0702_
timestamp 1676037725
transform -1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0703_
timestamp 1676037725
transform -1 0 17572 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0704_
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0705_
timestamp 1676037725
transform -1 0 16376 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 1676037725
transform -1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0708_
timestamp 1676037725
transform -1 0 14812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0709_
timestamp 1676037725
transform -1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0710_
timestamp 1676037725
transform 1 0 11960 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0713_
timestamp 1676037725
transform 1 0 12880 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0714_
timestamp 1676037725
transform 1 0 13524 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1676037725
transform -1 0 14352 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 1676037725
transform -1 0 13524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0717_
timestamp 1676037725
transform 1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0718_
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0719_
timestamp 1676037725
transform -1 0 13616 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0720_
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0721_
timestamp 1676037725
transform -1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0722_
timestamp 1676037725
transform -1 0 29256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1676037725
transform 1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29072 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1676037725
transform -1 0 28704 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1676037725
transform 1 0 24748 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0727_
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0728_
timestamp 1676037725
transform 1 0 25208 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0729_
timestamp 1676037725
transform 1 0 25668 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1676037725
transform 1 0 24932 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0731_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0732_
timestamp 1676037725
transform -1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1676037725
transform -1 0 28336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0734_
timestamp 1676037725
transform 1 0 28520 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30360 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0736_
timestamp 1676037725
transform -1 0 29072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0737_
timestamp 1676037725
transform 1 0 27416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1676037725
transform 1 0 27600 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0739_
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0740_
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 1676037725
transform -1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0742_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0743_
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0744_
timestamp 1676037725
transform 1 0 27508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0745_
timestamp 1676037725
transform 1 0 28152 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0746_
timestamp 1676037725
transform -1 0 26864 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0747_
timestamp 1676037725
transform 1 0 27140 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0748_
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp 1676037725
transform -1 0 24472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0750_
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0751_
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0752_
timestamp 1676037725
transform -1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0753_
timestamp 1676037725
transform -1 0 31372 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0754_
timestamp 1676037725
transform -1 0 30084 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0755_
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0756_
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0757_
timestamp 1676037725
transform 1 0 27600 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0758_
timestamp 1676037725
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1676037725
transform 1 0 28704 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0760_
timestamp 1676037725
transform -1 0 29256 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0761_
timestamp 1676037725
transform -1 0 26588 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 1676037725
transform 1 0 25760 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0763_
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0764_
timestamp 1676037725
transform 1 0 28888 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0765_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0766_
timestamp 1676037725
transform 1 0 30452 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0767_
timestamp 1676037725
transform -1 0 31372 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0768_
timestamp 1676037725
transform 1 0 30728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1676037725
transform 1 0 29808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0770_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0771_
timestamp 1676037725
transform -1 0 29440 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0772_
timestamp 1676037725
transform 1 0 29532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0773_
timestamp 1676037725
transform 1 0 29348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0774_
timestamp 1676037725
transform 1 0 24288 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0775_
timestamp 1676037725
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _0776_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0777_
timestamp 1676037725
transform -1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0778_
timestamp 1676037725
transform 1 0 27324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1676037725
transform -1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1676037725
transform -1 0 23368 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0782_
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0783_
timestamp 1676037725
transform 1 0 25668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1676037725
transform -1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0785_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0786_
timestamp 1676037725
transform 1 0 25576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0787_
timestamp 1676037725
transform -1 0 26220 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0788_
timestamp 1676037725
transform 1 0 25576 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0789_
timestamp 1676037725
transform -1 0 26312 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0790_
timestamp 1676037725
transform 1 0 20976 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0791_
timestamp 1676037725
transform -1 0 22632 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0792_
timestamp 1676037725
transform -1 0 23644 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0793_
timestamp 1676037725
transform -1 0 22632 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0794_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0795_
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0796_
timestamp 1676037725
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1676037725
transform -1 0 3496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0798_
timestamp 1676037725
transform -1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0799_
timestamp 1676037725
transform -1 0 2852 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 1676037725
transform -1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0801_
timestamp 1676037725
transform -1 0 9752 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1676037725
transform -1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0803_
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0804_
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0805_
timestamp 1676037725
transform 1 0 2392 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0806_
timestamp 1676037725
transform 1 0 2392 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0807_
timestamp 1676037725
transform -1 0 2852 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 1676037725
transform 1 0 2300 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0810_
timestamp 1676037725
transform 1 0 3312 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0811_
timestamp 1676037725
transform -1 0 8004 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0812_
timestamp 1676037725
transform 1 0 5612 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _0813_
timestamp 1676037725
transform -1 0 6716 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0814_
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1676037725
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0816_
timestamp 1676037725
transform -1 0 4416 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0817_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0818_
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0819_
timestamp 1676037725
transform -1 0 7084 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1676037725
transform 1 0 4784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0821_
timestamp 1676037725
transform -1 0 3496 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0822_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0824_
timestamp 1676037725
transform -1 0 3956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1676037725
transform -1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0826_
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0827_
timestamp 1676037725
transform 1 0 2668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0828_
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0829_
timestamp 1676037725
transform -1 0 6624 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 1676037725
transform 1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0831_
timestamp 1676037725
transform -1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0832_
timestamp 1676037725
transform -1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0833_
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0835_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0836_
timestamp 1676037725
transform -1 0 12604 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0837_
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1676037725
transform 1 0 16836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0839_
timestamp 1676037725
transform -1 0 24012 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1676037725
transform -1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1676037725
transform -1 0 24104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0842_
timestamp 1676037725
transform -1 0 23460 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0843_
timestamp 1676037725
transform -1 0 23184 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0844_
timestamp 1676037725
transform -1 0 21344 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0845_
timestamp 1676037725
transform 1 0 17020 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0846_
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0847_
timestamp 1676037725
transform -1 0 20884 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0848_
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0849_
timestamp 1676037725
transform -1 0 21068 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0850_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0851_
timestamp 1676037725
transform -1 0 20332 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0852_
timestamp 1676037725
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0853_
timestamp 1676037725
transform -1 0 17756 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0854_
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0856_
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0857_
timestamp 1676037725
transform 1 0 17480 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0858_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1676037725
transform -1 0 18952 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0860_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0861_
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0862_
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0863_
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0864_
timestamp 1676037725
transform -1 0 19136 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0865_
timestamp 1676037725
transform -1 0 16376 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0866_
timestamp 1676037725
transform -1 0 17112 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0867_
timestamp 1676037725
transform 1 0 13432 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0868_
timestamp 1676037725
transform -1 0 26680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0869_
timestamp 1676037725
transform -1 0 4692 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1676037725
transform -1 0 2852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0872_
timestamp 1676037725
transform -1 0 9568 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0873_
timestamp 1676037725
transform -1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1676037725
transform -1 0 7912 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1676037725
transform 1 0 6808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0876_
timestamp 1676037725
transform -1 0 7452 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 1676037725
transform -1 0 6164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1676037725
transform 1 0 7544 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0879_
timestamp 1676037725
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0880_
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1676037725
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0882_
timestamp 1676037725
transform -1 0 6072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0883_
timestamp 1676037725
transform -1 0 5336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1676037725
transform -1 0 2576 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0885_
timestamp 1676037725
transform 1 0 2760 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1676037725
transform 1 0 4232 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0888_
timestamp 1676037725
transform -1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0889_
timestamp 1676037725
transform -1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0891_
timestamp 1676037725
transform -1 0 2668 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0892_
timestamp 1676037725
transform -1 0 3404 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1676037725
transform -1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0894_
timestamp 1676037725
transform 1 0 2852 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0895_
timestamp 1676037725
transform -1 0 4508 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0896_
timestamp 1676037725
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0897_
timestamp 1676037725
transform -1 0 23920 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0898_
timestamp 1676037725
transform 1 0 21160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1676037725
transform 1 0 21988 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1676037725
transform -1 0 21528 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0902_
timestamp 1676037725
transform -1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0903_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0904_
timestamp 1676037725
transform -1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0905_
timestamp 1676037725
transform -1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0906_
timestamp 1676037725
transform -1 0 10856 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1676037725
transform -1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0908_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0910_
timestamp 1676037725
transform -1 0 10488 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1676037725
transform -1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0912_
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0914_
timestamp 1676037725
transform -1 0 11592 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1676037725
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0916_
timestamp 1676037725
transform -1 0 10672 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1676037725
transform -1 0 8280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0918_
timestamp 1676037725
transform -1 0 10764 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 1676037725
transform 1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0920_
timestamp 1676037725
transform 1 0 26680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0921_
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0922_
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0924_
timestamp 1676037725
transform -1 0 30636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1676037725
transform -1 0 24104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0926_
timestamp 1676037725
transform -1 0 29992 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0927_
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0928_
timestamp 1676037725
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0929_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0930_
timestamp 1676037725
transform -1 0 27600 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0931_
timestamp 1676037725
transform -1 0 28888 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0932_
timestamp 1676037725
transform 1 0 25024 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0933_
timestamp 1676037725
transform -1 0 25484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0934_
timestamp 1676037725
transform 1 0 26036 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0935_
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0936_
timestamp 1676037725
transform 1 0 23184 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0937_
timestamp 1676037725
transform 1 0 22448 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 1676037725
transform 1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_2  _0939_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _0940_
timestamp 1676037725
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0942_
timestamp 1676037725
transform -1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1676037725
transform -1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0944_
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0945_
timestamp 1676037725
transform -1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1676037725
transform -1 0 18032 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1676037725
transform -1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1676037725
transform 1 0 18400 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1676037725
transform 1 0 17572 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0950_
timestamp 1676037725
transform -1 0 16376 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0951_
timestamp 1676037725
transform -1 0 19964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0952_
timestamp 1676037725
transform -1 0 20056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0953_
timestamp 1676037725
transform -1 0 20884 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0955_
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0956_
timestamp 1676037725
transform -1 0 10856 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0957_
timestamp 1676037725
transform 1 0 12512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0958_
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0959_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0960_
timestamp 1676037725
transform -1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0961_
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0962_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1676037725
transform 1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0965_
timestamp 1676037725
transform -1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0966_
timestamp 1676037725
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0968_
timestamp 1676037725
transform -1 0 11040 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0969_
timestamp 1676037725
transform -1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0970_
timestamp 1676037725
transform -1 0 11132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1676037725
transform -1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0972_
timestamp 1676037725
transform -1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1676037725
transform -1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0974_
timestamp 1676037725
transform 1 0 8464 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 1676037725
transform 1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1676037725
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0977_
timestamp 1676037725
transform -1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1676037725
transform 1 0 9936 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0979_
timestamp 1676037725
transform -1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0980_
timestamp 1676037725
transform 1 0 9476 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0981_
timestamp 1676037725
transform -1 0 10488 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1676037725
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0983_
timestamp 1676037725
transform -1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0984_
timestamp 1676037725
transform -1 0 5336 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1676037725
transform -1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0986_
timestamp 1676037725
transform -1 0 8648 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0987_
timestamp 1676037725
transform 1 0 9108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0988_
timestamp 1676037725
transform 1 0 4692 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0989_
timestamp 1676037725
transform -1 0 6072 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0990_
timestamp 1676037725
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0991_
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _0992_
timestamp 1676037725
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0993_
timestamp 1676037725
transform 1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0994_
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0995_
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0997_
timestamp 1676037725
transform -1 0 4416 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0998_
timestamp 1676037725
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0999_
timestamp 1676037725
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1000_
timestamp 1676037725
transform -1 0 3496 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1001_
timestamp 1676037725
transform 1 0 3404 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1676037725
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1003_
timestamp 1676037725
transform 1 0 2392 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1004_
timestamp 1676037725
transform 1 0 7360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1676037725
transform -1 0 8832 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1676037725
transform -1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1007_
timestamp 1676037725
transform -1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1008_
timestamp 1676037725
transform -1 0 3036 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1009_
timestamp 1676037725
transform -1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1010_
timestamp 1676037725
transform -1 0 3496 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1011_
timestamp 1676037725
transform 1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1012_
timestamp 1676037725
transform -1 0 6992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1676037725
transform -1 0 6072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1014_
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1015_
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1016_
timestamp 1676037725
transform -1 0 3128 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1017_
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1018_
timestamp 1676037725
transform -1 0 3680 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 1676037725
transform -1 0 5980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1020_
timestamp 1676037725
transform -1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1676037725
transform -1 0 31372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1024_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform -1 0 23828 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform -1 0 21344 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1028_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1676037725
transform -1 0 16376 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 14444 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 11776 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1032_
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1033_
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1676037725
transform 1 0 22632 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1036_
timestamp 1676037725
transform 1 0 29532 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1037_
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1038_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1676037725
transform 1 0 27692 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1676037725
transform 1 0 6716 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1676037725
transform 1 0 14444 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1043_
timestamp 1676037725
transform -1 0 11224 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1046_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1047_
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1048_
timestamp 1676037725
transform -1 0 8280 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1049_
timestamp 1676037725
transform -1 0 7544 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 5888 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1051_
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1676037725
transform 1 0 4048 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1053_
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform -1 0 19780 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1057_
timestamp 1676037725
transform -1 0 11960 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1058_
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1059_
timestamp 1676037725
transform -1 0 10764 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1060_
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1676037725
transform -1 0 31188 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1676037725
transform -1 0 28888 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1676037725
transform 1 0 26496 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1676037725
transform 1 0 21988 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1068_
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1676037725
transform 1 0 19780 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1676037725
transform 1 0 11040 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1676037725
transform -1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1676037725
transform 1 0 7176 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1074_
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1676037725
transform -1 0 5980 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1076_
timestamp 1676037725
transform 1 0 4600 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1077_
timestamp 1676037725
transform 1 0 6900 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1078_
timestamp 1676037725
transform 1 0 6532 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1676037725
transform 1 0 4600 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1676037725
transform 1 0 15456 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1676037725
transform 1 0 14628 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1676037725
transform 1 0 30268 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1676037725
transform -1 0 31280 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1676037725
transform 1 0 29716 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1676037725
transform -1 0 31372 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1676037725
transform 1 0 29072 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1676037725
transform -1 0 29808 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1676037725
transform -1 0 31740 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1100_
timestamp 1676037725
transform -1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1676037725
transform -1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1102_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1103_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1104_
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1676037725
transform -1 0 16376 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1106_
timestamp 1676037725
transform -1 0 13800 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1108_
timestamp 1676037725
transform -1 0 13800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19780 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1676037725
transform -1 0 9660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1676037725
transform -1 0 9660 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1676037725
transform -1 0 22632 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1676037725
transform 1 0 23368 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1676037725
transform 1 0 28520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1676037725
transform 1 0 30912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform -1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform -1 0 31832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform -1 0 25944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform -1 0 29072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 28060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4324 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_8
timestamp 1676037725
transform -1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_9
timestamp 1676037725
transform -1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_10
timestamp 1676037725
transform -1 0 2208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_11
timestamp 1676037725
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_12
timestamp 1676037725
transform -1 0 2208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_13
timestamp 1676037725
transform -1 0 1840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_algofoogle_solo_squash_14
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 314 592
<< labels >>
flabel metal4 s 31710 21560 31770 21760 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 32446 21560 32506 21760 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30974 21560 31034 21760 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30238 21560 30298 21760 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 29502 21560 29562 21760 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 28766 21560 28826 21760 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 28030 21560 28090 21760 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 27294 21560 27354 21760 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 26558 21560 26618 21760 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 25822 21560 25882 21760 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 25086 21560 25146 21760 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 24350 21560 24410 21760 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 23614 21560 23674 21760 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22878 21560 22938 21760 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 22142 21560 22202 21760 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21406 21560 21466 21760 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20670 21560 20730 21760 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 21560 19994 21760 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19198 21560 19258 21760 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 6686 21560 6746 21760 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 5950 21560 6010 21760 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 5214 21560 5274 21760 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 4478 21560 4538 21760 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 3742 21560 3802 21760 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 3006 21560 3066 21760 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 2270 21560 2330 21760 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 1534 21560 1594 21760 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 12574 21560 12634 21760 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 11838 21560 11898 21760 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 11102 21560 11162 21760 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 10366 21560 10426 21760 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 9630 21560 9690 21760 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 8894 21560 8954 21760 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 8158 21560 8218 21760 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 7422 21560 7482 21760 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 18462 21560 18522 21760 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 17726 21560 17786 21760 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 16990 21560 17050 21760 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 16254 21560 16314 21760 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 15518 21560 15578 21760 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 14782 21560 14842 21760 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 14046 21560 14106 21760 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 13310 21560 13370 21760 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 s 4865 1040 5185 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 12707 1040 13027 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 20549 1040 20869 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 28391 1040 28711 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8786 1040 9106 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 16628 1040 16948 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 24470 1040 24790 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 32312 1040 32632 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
rlabel metal1 16790 20128 16790 20128 0 vccd1
rlabel via1 16868 20672 16868 20672 0 vssd1
rlabel via1 22489 8942 22489 8942 0 _0000_
rlabel metal1 24058 7990 24058 7990 0 _0001_
rlabel metal2 21206 8262 21206 8262 0 _0002_
rlabel metal2 19918 8466 19918 8466 0 _0003_
rlabel metal1 17572 8058 17572 8058 0 _0004_
rlabel metal1 16156 8466 16156 8466 0 _0005_
rlabel metal1 14664 7854 14664 7854 0 _0006_
rlabel metal1 11668 7786 11668 7786 0 _0007_
rlabel metal2 25438 8262 25438 8262 0 _0008_
rlabel metal1 27140 8058 27140 8058 0 _0009_
rlabel metal2 24334 9078 24334 9078 0 _0010_
rlabel metal1 30723 9622 30723 9622 0 _0011_
rlabel metal1 30125 8466 30125 8466 0 _0012_
rlabel via1 30585 12818 30585 12818 0 _0013_
rlabel metal1 29936 14382 29936 14382 0 _0014_
rlabel metal2 27830 13702 27830 13702 0 _0015_
rlabel via1 13473 12818 13473 12818 0 _0016_
rlabel via1 7033 12818 7033 12818 0 _0017_
rlabel via1 14761 8942 14761 8942 0 _0018_
rlabel metal2 12558 11934 12558 11934 0 _0019_
rlabel via1 13289 9554 13289 9554 0 _0020_
rlabel metal1 3618 19414 3618 19414 0 _0021_
rlabel metal1 9328 19822 9328 19822 0 _0022_
rlabel metal1 6746 19754 6746 19754 0 _0023_
rlabel metal1 8786 18122 8786 18122 0 _0024_
rlabel metal2 8418 14994 8418 14994 0 _0025_
rlabel metal2 5290 16218 5290 16218 0 _0026_
rlabel metal2 4278 16354 4278 16354 0 _0027_
rlabel metal1 2346 16626 2346 16626 0 _0028_
rlabel metal2 3542 19618 3542 19618 0 _0029_
rlabel metal2 4462 18054 4462 18054 0 _0030_
rlabel via1 19462 12886 19462 12886 0 _0031_
rlabel metal1 9420 13906 9420 13906 0 _0032_
rlabel metal1 11684 14042 11684 14042 0 _0033_
rlabel metal1 8781 17238 8781 17238 0 _0034_
rlabel metal1 8418 15130 8418 15130 0 _0035_
rlabel metal2 10442 11730 10442 11730 0 _0036_
rlabel metal1 29936 16558 29936 16558 0 _0037_
rlabel metal2 31050 15878 31050 15878 0 _0038_
rlabel metal2 28290 16932 28290 16932 0 _0039_
rlabel metal2 26634 17442 26634 17442 0 _0040_
rlabel via1 23409 17238 23409 17238 0 _0041_
rlabel metal2 22126 16762 22126 16762 0 _0042_
rlabel metal1 14480 14382 14480 14382 0 _0043_
rlabel metal1 17608 13294 17608 13294 0 _0044_
rlabel metal1 16734 14382 16734 14382 0 _0045_
rlabel metal1 20235 14382 20235 14382 0 _0046_
rlabel metal1 11086 9486 11086 9486 0 _0047_
rlabel via1 11826 8942 11826 8942 0 _0048_
rlabel metal1 6946 7514 6946 7514 0 _0049_
rlabel metal1 9000 9962 9000 9962 0 _0050_
rlabel metal1 6486 6970 6486 6970 0 _0051_
rlabel metal1 5101 9962 5101 9962 0 _0052_
rlabel metal1 6900 8058 6900 8058 0 _0053_
rlabel via1 6849 9962 6849 9962 0 _0054_
rlabel metal1 4830 11322 4830 11322 0 _0055_
rlabel metal1 31326 13804 31326 13804 0 _0056_
rlabel metal1 14904 13702 14904 13702 0 _0057_
rlabel metal2 13202 15130 13202 15130 0 _0058_
rlabel metal2 13754 17306 13754 17306 0 _0059_
rlabel metal1 15594 16966 15594 16966 0 _0060_
rlabel metal2 14766 17510 14766 17510 0 _0061_
rlabel metal1 10212 19346 10212 19346 0 _0062_
rlabel metal1 8970 18938 8970 18938 0 _0063_
rlabel metal1 8740 18734 8740 18734 0 _0064_
rlabel metal2 9982 18462 9982 18462 0 _0065_
rlabel metal2 10074 17952 10074 17952 0 _0066_
rlabel metal1 18722 17000 18722 17000 0 _0067_
rlabel metal1 21482 19380 21482 19380 0 _0068_
rlabel metal2 20930 18054 20930 18054 0 _0069_
rlabel metal1 10304 20298 10304 20298 0 _0070_
rlabel metal1 12374 19380 12374 19380 0 _0071_
rlabel metal2 14214 16252 14214 16252 0 _0072_
rlabel metal2 11454 18054 11454 18054 0 _0073_
rlabel metal1 12696 18394 12696 18394 0 _0074_
rlabel via2 13386 18717 13386 18717 0 _0075_
rlabel metal1 10626 17748 10626 17748 0 _0076_
rlabel metal1 13478 18700 13478 18700 0 _0077_
rlabel metal2 12558 17731 12558 17731 0 _0078_
rlabel metal1 15916 16150 15916 16150 0 _0079_
rlabel metal1 16146 14246 16146 14246 0 _0080_
rlabel metal1 13340 16558 13340 16558 0 _0081_
rlabel metal1 13892 16218 13892 16218 0 _0082_
rlabel metal1 2622 12308 2622 12308 0 _0083_
rlabel viali 13758 17170 13758 17170 0 _0084_
rlabel metal1 2392 17578 2392 17578 0 _0085_
rlabel metal1 13573 17306 13573 17306 0 _0086_
rlabel metal1 21390 9622 21390 9622 0 _0087_
rlabel metal1 19918 15946 19918 15946 0 _0088_
rlabel metal1 18814 17102 18814 17102 0 _0089_
rlabel metal2 21022 15674 21022 15674 0 _0090_
rlabel metal1 17756 17306 17756 17306 0 _0091_
rlabel metal1 7682 19312 7682 19312 0 _0092_
rlabel metal2 16330 18122 16330 18122 0 _0093_
rlabel metal1 7544 17782 7544 17782 0 _0094_
rlabel viali 15778 18258 15778 18258 0 _0095_
rlabel metal1 19274 17680 19274 17680 0 _0096_
rlabel metal1 16238 17136 16238 17136 0 _0097_
rlabel metal1 16146 17306 16146 17306 0 _0098_
rlabel metal2 12742 17408 12742 17408 0 _0099_
rlabel metal2 12926 17442 12926 17442 0 _0100_
rlabel metal1 12512 16762 12512 16762 0 _0101_
rlabel viali 15226 17647 15226 17647 0 _0102_
rlabel viali 12374 17638 12374 17638 0 _0103_
rlabel metal1 12098 17850 12098 17850 0 _0104_
rlabel metal1 14168 15470 14168 15470 0 _0105_
rlabel metal2 15134 16150 15134 16150 0 _0106_
rlabel metal1 20746 16048 20746 16048 0 _0107_
rlabel metal1 19149 16218 19149 16218 0 _0108_
rlabel metal1 17480 17646 17480 17646 0 _0109_
rlabel metal1 17250 17612 17250 17612 0 _0110_
rlabel metal2 17710 17340 17710 17340 0 _0111_
rlabel metal2 20010 17374 20010 17374 0 _0112_
rlabel metal1 17526 16082 17526 16082 0 _0113_
rlabel metal1 14490 14042 14490 14042 0 _0114_
rlabel metal1 15410 14824 15410 14824 0 _0115_
rlabel metal1 9591 16558 9591 16558 0 _0116_
rlabel metal1 15318 15028 15318 15028 0 _0117_
rlabel metal1 14904 13158 14904 13158 0 _0118_
rlabel metal1 15916 14790 15916 14790 0 _0119_
rlabel metal1 16284 16218 16284 16218 0 _0120_
rlabel metal2 16514 16116 16514 16116 0 _0121_
rlabel metal1 14812 18802 14812 18802 0 _0122_
rlabel metal1 25852 19346 25852 19346 0 _0123_
rlabel metal2 20930 18547 20930 18547 0 _0124_
rlabel metal1 24012 18394 24012 18394 0 _0125_
rlabel metal2 20286 17476 20286 17476 0 _0126_
rlabel metal1 19550 17748 19550 17748 0 _0127_
rlabel metal1 23276 18734 23276 18734 0 _0128_
rlabel metal1 24150 18666 24150 18666 0 _0129_
rlabel metal1 23460 20434 23460 20434 0 _0130_
rlabel metal2 25898 19567 25898 19567 0 _0131_
rlabel metal2 23046 20060 23046 20060 0 _0132_
rlabel metal2 22126 18870 22126 18870 0 _0133_
rlabel metal1 22264 19822 22264 19822 0 _0134_
rlabel metal1 20194 19482 20194 19482 0 _0135_
rlabel metal1 20516 18394 20516 18394 0 _0136_
rlabel metal1 20562 19346 20562 19346 0 _0137_
rlabel metal2 21206 19108 21206 19108 0 _0138_
rlabel metal2 22770 18836 22770 18836 0 _0139_
rlabel metal2 22034 18938 22034 18938 0 _0140_
rlabel metal2 19826 18088 19826 18088 0 _0141_
rlabel metal2 22402 19380 22402 19380 0 _0142_
rlabel metal1 21850 19686 21850 19686 0 _0143_
rlabel metal2 18722 19380 18722 19380 0 _0144_
rlabel metal1 20010 19992 20010 19992 0 _0145_
rlabel metal2 18906 19516 18906 19516 0 _0146_
rlabel metal1 19550 18938 19550 18938 0 _0147_
rlabel metal1 20148 20502 20148 20502 0 _0148_
rlabel metal2 22126 20196 22126 20196 0 _0149_
rlabel metal2 24978 20026 24978 20026 0 _0150_
rlabel metal1 23138 19244 23138 19244 0 _0151_
rlabel metal1 23598 19278 23598 19278 0 _0152_
rlabel metal1 26082 19482 26082 19482 0 _0153_
rlabel metal2 26542 19142 26542 19142 0 _0154_
rlabel metal2 26450 18836 26450 18836 0 _0155_
rlabel metal1 27002 19482 27002 19482 0 _0156_
rlabel metal1 25162 19278 25162 19278 0 _0157_
rlabel metal1 24748 19210 24748 19210 0 _0158_
rlabel metal1 21114 19890 21114 19890 0 _0159_
rlabel metal2 20194 20230 20194 20230 0 _0160_
rlabel metal1 14950 19992 14950 19992 0 _0161_
rlabel metal1 20562 20026 20562 20026 0 _0162_
rlabel metal1 10074 20298 10074 20298 0 _0163_
rlabel metal1 16698 18768 16698 18768 0 _0164_
rlabel metal1 20378 16150 20378 16150 0 _0165_
rlabel metal2 19734 16388 19734 16388 0 _0166_
rlabel metal2 2254 18326 2254 18326 0 _0167_
rlabel metal1 2530 17068 2530 17068 0 _0168_
rlabel metal1 3036 17850 3036 17850 0 _0169_
rlabel metal1 3496 18394 3496 18394 0 _0170_
rlabel metal1 17710 9996 17710 9996 0 _0171_
rlabel metal1 15410 10166 15410 10166 0 _0172_
rlabel metal1 14812 10234 14812 10234 0 _0173_
rlabel metal2 2898 7548 2898 7548 0 _0174_
rlabel metal1 6624 11254 6624 11254 0 _0175_
rlabel metal2 15318 11050 15318 11050 0 _0176_
rlabel metal2 15870 11288 15870 11288 0 _0177_
rlabel metal2 2714 16898 2714 16898 0 _0178_
rlabel metal1 12834 14994 12834 14994 0 _0179_
rlabel metal1 23414 14382 23414 14382 0 _0180_
rlabel metal1 24978 15946 24978 15946 0 _0181_
rlabel metal1 24564 14586 24564 14586 0 _0182_
rlabel metal1 24610 14382 24610 14382 0 _0183_
rlabel metal1 24288 13702 24288 13702 0 _0184_
rlabel metal1 12972 13294 12972 13294 0 _0185_
rlabel metal1 10012 13226 10012 13226 0 _0186_
rlabel metal2 13570 10013 13570 10013 0 _0187_
rlabel metal1 14536 11526 14536 11526 0 _0188_
rlabel metal1 16928 7854 16928 7854 0 _0189_
rlabel metal2 22218 10166 22218 10166 0 _0190_
rlabel metal1 17986 15504 17986 15504 0 _0191_
rlabel metal2 21298 15351 21298 15351 0 _0192_
rlabel via2 7774 17595 7774 17595 0 _0193_
rlabel metal2 14766 13498 14766 13498 0 _0194_
rlabel metal1 14858 9554 14858 9554 0 _0195_
rlabel metal1 5290 9622 5290 9622 0 _0196_
rlabel metal1 13938 7412 13938 7412 0 _0197_
rlabel metal1 23322 7514 23322 7514 0 _0198_
rlabel metal1 24748 7378 24748 7378 0 _0199_
rlabel metal2 24334 7786 24334 7786 0 _0200_
rlabel metal1 24050 7718 24050 7718 0 _0201_
rlabel metal1 23046 7752 23046 7752 0 _0202_
rlabel metal1 23828 7854 23828 7854 0 _0203_
rlabel metal1 14812 6834 14812 6834 0 _0204_
rlabel metal1 21574 6800 21574 6800 0 _0205_
rlabel metal1 21482 5270 21482 5270 0 _0206_
rlabel metal2 21758 6970 21758 6970 0 _0207_
rlabel metal1 22011 6834 22011 6834 0 _0208_
rlabel metal1 21712 5678 21712 5678 0 _0209_
rlabel metal2 22402 7344 22402 7344 0 _0210_
rlabel metal1 20976 7854 20976 7854 0 _0211_
rlabel metal2 19458 8364 19458 8364 0 _0212_
rlabel metal1 25576 13906 25576 13906 0 _0213_
rlabel metal2 22678 14042 22678 14042 0 _0214_
rlabel metal2 22494 14586 22494 14586 0 _0215_
rlabel metal1 20378 7378 20378 7378 0 _0216_
rlabel metal1 20884 5882 20884 5882 0 _0217_
rlabel metal1 21068 6766 21068 6766 0 _0218_
rlabel metal2 20470 7072 20470 7072 0 _0219_
rlabel metal2 21666 6698 21666 6698 0 _0220_
rlabel metal1 19780 7514 19780 7514 0 _0221_
rlabel metal1 17756 6222 17756 6222 0 _0222_
rlabel metal2 17158 6052 17158 6052 0 _0223_
rlabel metal2 17066 6052 17066 6052 0 _0224_
rlabel metal1 20792 5338 20792 5338 0 _0225_
rlabel metal2 21206 6732 21206 6732 0 _0226_
rlabel metal1 17664 6290 17664 6290 0 _0227_
rlabel metal1 17342 6970 17342 6970 0 _0228_
rlabel metal2 17894 7684 17894 7684 0 _0229_
rlabel metal1 16974 5678 16974 5678 0 _0230_
rlabel metal1 18078 6732 18078 6732 0 _0231_
rlabel metal1 16146 7310 16146 7310 0 _0232_
rlabel metal1 16560 7174 16560 7174 0 _0233_
rlabel metal2 15410 7650 15410 7650 0 _0234_
rlabel metal1 16376 7514 16376 7514 0 _0235_
rlabel metal1 17020 8058 17020 8058 0 _0236_
rlabel metal2 12466 6732 12466 6732 0 _0237_
rlabel metal2 12006 6460 12006 6460 0 _0238_
rlabel metal1 12788 6290 12788 6290 0 _0239_
rlabel metal2 16238 5916 16238 5916 0 _0240_
rlabel metal2 13202 6052 13202 6052 0 _0241_
rlabel metal1 13616 6426 13616 6426 0 _0242_
rlabel metal2 14122 7990 14122 7990 0 _0243_
rlabel metal1 13616 8466 13616 8466 0 _0244_
rlabel metal1 12903 6766 12903 6766 0 _0245_
rlabel metal1 12926 6834 12926 6834 0 _0246_
rlabel metal2 13110 7140 13110 7140 0 _0247_
rlabel metal1 11776 7514 11776 7514 0 _0248_
rlabel metal1 29624 13430 29624 13430 0 _0249_
rlabel metal1 31924 18598 31924 18598 0 _0250_
rlabel metal1 28888 12818 28888 12818 0 _0251_
rlabel metal2 25254 13430 25254 13430 0 _0252_
rlabel metal2 25346 10846 25346 10846 0 _0253_
rlabel metal2 25162 14824 25162 14824 0 _0254_
rlabel metal2 31970 10642 31970 10642 0 _0255_
rlabel metal1 26128 10030 26128 10030 0 _0256_
rlabel metal2 24794 9146 24794 9146 0 _0257_
rlabel metal2 25254 8330 25254 8330 0 _0258_
rlabel metal1 17066 11016 17066 11016 0 _0259_
rlabel metal1 27324 12818 27324 12818 0 _0260_
rlabel metal1 29854 13362 29854 13362 0 _0261_
rlabel metal1 27922 9010 27922 9010 0 _0262_
rlabel metal1 28106 8058 28106 8058 0 _0263_
rlabel metal1 26818 9010 26818 9010 0 _0264_
rlabel metal2 26634 9384 26634 9384 0 _0265_
rlabel metal2 26818 8602 26818 8602 0 _0266_
rlabel metal1 27462 10642 27462 10642 0 _0267_
rlabel metal2 27922 10166 27922 10166 0 _0268_
rlabel metal2 27646 10336 27646 10336 0 _0269_
rlabel metal1 28980 9894 28980 9894 0 _0270_
rlabel metal2 27462 10642 27462 10642 0 _0271_
rlabel metal1 26358 10098 26358 10098 0 _0272_
rlabel metal1 24656 8466 24656 8466 0 _0273_
rlabel metal1 31786 9996 31786 9996 0 _0274_
rlabel metal2 31786 10438 31786 10438 0 _0275_
rlabel metal2 31050 10336 31050 10336 0 _0276_
rlabel metal2 29670 9724 29670 9724 0 _0277_
rlabel metal2 29762 9146 29762 9146 0 _0278_
rlabel metal2 29026 9860 29026 9860 0 _0279_
rlabel metal1 29532 11254 29532 11254 0 _0280_
rlabel metal1 28934 11084 28934 11084 0 _0281_
rlabel metal2 28750 10812 28750 10812 0 _0282_
rlabel metal2 26358 10268 26358 10268 0 _0283_
rlabel metal2 25990 9418 25990 9418 0 _0284_
rlabel metal1 30590 8908 30590 8908 0 _0285_
rlabel via1 29029 12070 29029 12070 0 _0286_
rlabel metal2 30222 11492 30222 11492 0 _0287_
rlabel metal2 31050 11356 31050 11356 0 _0288_
rlabel metal2 30774 11764 30774 11764 0 _0289_
rlabel metal1 30084 11866 30084 11866 0 _0290_
rlabel metal1 28750 11764 28750 11764 0 _0291_
rlabel metal1 29486 13906 29486 13906 0 _0292_
rlabel metal1 29578 13804 29578 13804 0 _0293_
rlabel metal1 24196 12954 24196 12954 0 _0294_
rlabel metal2 28198 11968 28198 11968 0 _0295_
rlabel metal1 27692 12818 27692 12818 0 _0296_
rlabel metal2 27646 12988 27646 12988 0 _0297_
rlabel metal2 29026 14450 29026 14450 0 _0298_
rlabel metal1 25760 12886 25760 12886 0 _0299_
rlabel metal1 23046 13906 23046 13906 0 _0300_
rlabel metal2 25714 13804 25714 13804 0 _0301_
rlabel metal1 26266 12954 26266 12954 0 _0302_
rlabel via2 25990 14331 25990 14331 0 _0303_
rlabel metal1 25392 14382 25392 14382 0 _0304_
rlabel metal1 26128 13362 26128 13362 0 _0305_
rlabel metal2 25622 11492 25622 11492 0 _0306_
rlabel metal1 26312 12410 26312 12410 0 _0307_
rlabel metal1 22448 13294 22448 13294 0 _0308_
rlabel metal1 21528 13294 21528 13294 0 _0309_
rlabel metal1 22448 13362 22448 13362 0 _0310_
rlabel metal1 22586 13192 22586 13192 0 _0311_
rlabel metal1 19596 13158 19596 13158 0 _0312_
rlabel metal1 14490 12818 14490 12818 0 _0313_
rlabel metal2 13754 12852 13754 12852 0 _0314_
rlabel metal1 1794 13872 1794 13872 0 _0315_
rlabel metal2 2254 13260 2254 13260 0 _0316_
rlabel metal2 2438 13260 2438 13260 0 _0317_
rlabel metal1 2553 12886 2553 12886 0 _0318_
rlabel metal2 9338 13056 9338 13056 0 _0319_
rlabel metal2 9798 12308 9798 12308 0 _0320_
rlabel metal1 9614 13294 9614 13294 0 _0321_
rlabel metal1 6440 13158 6440 13158 0 _0322_
rlabel metal1 3680 13226 3680 13226 0 _0323_
rlabel metal2 3450 14076 3450 14076 0 _0324_
rlabel metal1 2208 13294 2208 13294 0 _0325_
rlabel metal1 6118 13396 6118 13396 0 _0326_
rlabel metal2 5658 14416 5658 14416 0 _0327_
rlabel metal2 4554 14348 4554 14348 0 _0328_
rlabel metal2 6762 14008 6762 14008 0 _0329_
rlabel metal2 6026 13532 6026 13532 0 _0330_
rlabel metal1 6624 12138 6624 12138 0 _0331_
rlabel metal2 7130 13940 7130 13940 0 _0332_
rlabel metal1 6440 14518 6440 14518 0 _0333_
rlabel metal1 3266 13940 3266 13940 0 _0334_
rlabel metal2 4462 14042 4462 14042 0 _0335_
rlabel metal2 5382 13498 5382 13498 0 _0336_
rlabel metal1 6164 12886 6164 12886 0 _0337_
rlabel metal1 3174 12886 3174 12886 0 _0338_
rlabel metal1 3588 11866 3588 11866 0 _0339_
rlabel metal1 4922 12410 4922 12410 0 _0340_
rlabel metal1 5658 13498 5658 13498 0 _0341_
rlabel metal1 4738 13362 4738 13362 0 _0342_
rlabel metal2 3266 12988 3266 12988 0 _0343_
rlabel metal2 2714 13124 2714 13124 0 _0344_
rlabel metal1 4554 13294 4554 13294 0 _0345_
rlabel metal1 5980 12274 5980 12274 0 _0346_
rlabel metal1 6716 12206 6716 12206 0 _0347_
rlabel metal2 15226 10574 15226 10574 0 _0348_
rlabel metal1 15410 9554 15410 9554 0 _0349_
rlabel metal2 12098 12682 12098 12682 0 _0350_
rlabel metal1 13984 13158 13984 13158 0 _0351_
rlabel metal1 16882 15504 16882 15504 0 _0352_
rlabel metal1 19550 15504 19550 15504 0 _0353_
rlabel metal1 22862 11152 22862 11152 0 _0354_
rlabel metal2 22770 11322 22770 11322 0 _0355_
rlabel metal1 23828 10234 23828 10234 0 _0356_
rlabel metal1 23092 10234 23092 10234 0 _0357_
rlabel metal2 19090 11390 19090 11390 0 _0358_
rlabel metal2 20194 10744 20194 10744 0 _0359_
rlabel metal2 17802 11900 17802 11900 0 _0360_
rlabel metal1 17066 10574 17066 10574 0 _0361_
rlabel metal1 20010 10030 20010 10030 0 _0362_
rlabel metal1 18157 9894 18157 9894 0 _0363_
rlabel metal2 19826 9792 19826 9792 0 _0364_
rlabel metal1 19826 10234 19826 10234 0 _0365_
rlabel metal2 19458 11764 19458 11764 0 _0366_
rlabel metal1 16974 11322 16974 11322 0 _0367_
rlabel metal2 17342 9724 17342 9724 0 _0368_
rlabel metal2 16882 11628 16882 11628 0 _0369_
rlabel metal1 17572 11798 17572 11798 0 _0370_
rlabel metal1 17480 11322 17480 11322 0 _0371_
rlabel metal1 16330 11560 16330 11560 0 _0372_
rlabel metal1 17710 10778 17710 10778 0 _0373_
rlabel metal2 18538 10404 18538 10404 0 _0374_
rlabel metal1 18860 9486 18860 9486 0 _0375_
rlabel metal1 18998 9622 18998 9622 0 _0376_
rlabel metal1 18906 10642 18906 10642 0 _0377_
rlabel metal1 18584 10778 18584 10778 0 _0378_
rlabel metal1 16560 11730 16560 11730 0 _0379_
rlabel metal1 16406 11050 16406 11050 0 _0380_
rlabel metal1 15180 11254 15180 11254 0 _0381_
rlabel metal1 9276 19414 9276 19414 0 _0382_
rlabel metal1 2691 19822 2691 19822 0 _0383_
rlabel metal2 6854 19788 6854 19788 0 _0384_
rlabel metal1 7866 19482 7866 19482 0 _0385_
rlabel metal2 7222 18598 7222 18598 0 _0386_
rlabel metal1 7071 18394 7071 18394 0 _0387_
rlabel metal2 7038 18972 7038 18972 0 _0388_
rlabel metal1 8188 17646 8188 17646 0 _0389_
rlabel metal1 8280 14382 8280 14382 0 _0390_
rlabel metal1 5520 16150 5520 16150 0 _0391_
rlabel metal2 2070 16320 2070 16320 0 _0392_
rlabel metal2 2898 16320 2898 16320 0 _0393_
rlabel metal1 4186 16082 4186 16082 0 _0394_
rlabel metal2 2346 16320 2346 16320 0 _0395_
rlabel metal1 3404 18734 3404 18734 0 _0396_
rlabel metal2 2622 18666 2622 18666 0 _0397_
rlabel metal2 2254 19108 2254 19108 0 _0398_
rlabel viali 4202 17646 4202 17646 0 _0399_
rlabel metal2 23230 12580 23230 12580 0 _0400_
rlabel metal1 23184 12682 23184 12682 0 _0401_
rlabel metal1 21850 12682 21850 12682 0 _0402_
rlabel metal1 22448 12410 22448 12410 0 _0403_
rlabel metal2 21390 12988 21390 12988 0 _0404_
rlabel metal1 21206 12954 21206 12954 0 _0405_
rlabel metal1 19964 13294 19964 13294 0 _0406_
rlabel metal1 9200 15062 9200 15062 0 _0407_
rlabel metal1 10212 17238 10212 17238 0 _0408_
rlabel metal2 9982 14824 9982 14824 0 _0409_
rlabel metal1 11316 13906 11316 13906 0 _0410_
rlabel metal1 9246 16762 9246 16762 0 _0411_
rlabel metal2 9798 16966 9798 16966 0 _0412_
rlabel metal1 8970 16694 8970 16694 0 _0413_
rlabel metal1 10902 15334 10902 15334 0 _0414_
rlabel metal1 10626 16218 10626 16218 0 _0415_
rlabel metal1 8280 14994 8280 14994 0 _0416_
rlabel metal1 10350 11118 10350 11118 0 _0417_
rlabel metal1 27554 14586 27554 14586 0 _0418_
rlabel metal1 29134 15062 29134 15062 0 _0419_
rlabel metal1 28566 15130 28566 15130 0 _0420_
rlabel metal1 28382 16014 28382 16014 0 _0421_
rlabel metal1 23414 15572 23414 15572 0 _0422_
rlabel metal1 29256 15402 29256 15402 0 _0423_
rlabel metal1 28842 15572 28842 15572 0 _0424_
rlabel metal1 28198 16218 28198 16218 0 _0425_
rlabel metal1 26726 15130 26726 15130 0 _0426_
rlabel metal2 25070 15878 25070 15878 0 _0427_
rlabel metal1 25530 16218 25530 16218 0 _0428_
rlabel metal2 21114 15776 21114 15776 0 _0429_
rlabel metal2 23230 15912 23230 15912 0 _0430_
rlabel metal1 23552 16218 23552 16218 0 _0431_
rlabel metal1 17434 14994 17434 14994 0 _0432_
rlabel metal1 21298 15674 21298 15674 0 _0433_
rlabel metal1 13018 14042 13018 14042 0 _0434_
rlabel metal2 18538 15402 18538 15402 0 _0435_
rlabel metal1 17434 15130 17434 15130 0 _0436_
rlabel metal2 17342 14620 17342 14620 0 _0437_
rlabel metal1 19366 15470 19366 15470 0 _0438_
rlabel metal1 16974 15062 16974 15062 0 _0439_
rlabel metal1 20470 14790 20470 14790 0 _0440_
rlabel metal1 20086 15062 20086 15062 0 _0441_
rlabel metal1 20470 14926 20470 14926 0 _0442_
rlabel metal1 10120 8602 10120 8602 0 _0443_
rlabel metal2 12558 9724 12558 9724 0 _0444_
rlabel metal1 13110 9146 13110 9146 0 _0445_
rlabel metal1 9522 9384 9522 9384 0 _0446_
rlabel metal2 12926 9758 12926 9758 0 _0447_
rlabel metal1 11684 8534 11684 8534 0 _0448_
rlabel metal2 11730 9486 11730 9486 0 _0449_
rlabel metal2 7682 7650 7682 7650 0 _0450_
rlabel metal1 2254 7412 2254 7412 0 _0451_
rlabel metal2 9154 8296 9154 8296 0 _0452_
rlabel metal1 9062 7344 9062 7344 0 _0453_
rlabel metal1 11040 7446 11040 7446 0 _0454_
rlabel metal2 9522 7786 9522 7786 0 _0455_
rlabel metal1 10166 7208 10166 7208 0 _0456_
rlabel metal1 8188 7446 8188 7446 0 _0457_
rlabel metal1 6946 7344 6946 7344 0 _0458_
rlabel metal2 9522 6528 9522 6528 0 _0459_
rlabel metal1 9338 6324 9338 6324 0 _0460_
rlabel via1 10174 7446 10174 7446 0 _0461_
rlabel metal2 10258 7378 10258 7378 0 _0462_
rlabel metal2 10442 6970 10442 6970 0 _0463_
rlabel metal1 10028 6834 10028 6834 0 _0464_
rlabel metal1 10166 9146 10166 9146 0 _0465_
rlabel metal2 10074 10914 10074 10914 0 _0466_
rlabel metal1 2553 7174 2553 7174 0 _0467_
rlabel metal1 4646 6358 4646 6358 0 _0468_
rlabel metal1 4232 6970 4232 6970 0 _0469_
rlabel metal1 8970 6834 8970 6834 0 _0470_
rlabel metal1 5520 6834 5520 6834 0 _0471_
rlabel metal1 5336 6970 5336 6970 0 _0472_
rlabel metal2 6578 6970 6578 6970 0 _0473_
rlabel metal1 3588 7514 3588 7514 0 _0474_
rlabel metal1 4232 6426 4232 6426 0 _0475_
rlabel metal1 5060 7514 5060 7514 0 _0476_
rlabel metal2 5474 8738 5474 8738 0 _0477_
rlabel metal1 5796 9146 5796 9146 0 _0478_
rlabel metal2 3266 8398 3266 8398 0 _0479_
rlabel metal2 2898 8908 2898 8908 0 _0480_
rlabel metal2 2254 9248 2254 9248 0 _0481_
rlabel metal1 1794 8398 1794 8398 0 _0482_
rlabel metal1 2024 8466 2024 8466 0 _0483_
rlabel metal1 2208 8398 2208 8398 0 _0484_
rlabel metal1 3036 8602 3036 8602 0 _0485_
rlabel metal1 8280 8466 8280 8466 0 _0486_
rlabel metal1 6854 7854 6854 7854 0 _0487_
rlabel metal2 3174 9214 3174 9214 0 _0488_
rlabel metal1 2438 9656 2438 9656 0 _0489_
rlabel metal1 3910 9622 3910 9622 0 _0490_
rlabel metal1 3818 9146 3818 9146 0 _0491_
rlabel metal1 5750 8942 5750 8942 0 _0492_
rlabel metal1 6532 9146 6532 9146 0 _0493_
rlabel metal2 2346 10166 2346 10166 0 _0494_
rlabel metal2 2714 10370 2714 10370 0 _0495_
rlabel metal2 2622 10778 2622 10778 0 _0496_
rlabel metal2 3450 10880 3450 10880 0 _0497_
rlabel metal1 3818 10778 3818 10778 0 _0498_
rlabel metal1 4922 11050 4922 11050 0 _0499_
rlabel metal1 4600 11118 4600 11118 0 _0500_
rlabel metal1 30912 13906 30912 13906 0 _0501_
rlabel metal2 31786 15963 31786 15963 0 clk
rlabel metal3 15778 13940 15778 13940 0 clknet_0_clk
rlabel metal1 6670 12750 6670 12750 0 clknet_3_0__leaf_clk
rlabel metal1 13018 9588 13018 9588 0 clknet_3_1__leaf_clk
rlabel metal1 8786 15878 8786 15878 0 clknet_3_2__leaf_clk
rlabel metal1 16422 19822 16422 19822 0 clknet_3_3__leaf_clk
rlabel metal1 20332 12750 20332 12750 0 clknet_3_4__leaf_clk
rlabel metal1 29578 8500 29578 8500 0 clknet_3_5__leaf_clk
rlabel metal1 27646 15334 27646 15334 0 clknet_3_6__leaf_clk
rlabel metal1 22034 16694 22034 16694 0 clknet_3_7__leaf_clk
rlabel metal1 30539 18326 30539 18326 0 down_key.d
rlabel metal1 30958 18156 30958 18156 0 down_key.dff1
rlabel metal1 29992 13294 29992 13294 0 down_key.dff2
rlabel metal2 12466 11798 12466 11798 0 game.ballDirX
rlabel metal2 17618 7378 17618 7378 0 game.ballDirY
rlabel metal1 12466 9962 12466 9962 0 game.ballX\[0\]
rlabel metal1 12558 8500 12558 8500 0 game.ballX\[1\]
rlabel metal1 8096 14450 8096 14450 0 game.ballX\[2\]
rlabel metal1 10350 10234 10350 10234 0 game.ballX\[3\]
rlabel metal2 5290 7038 5290 7038 0 game.ballX\[4\]
rlabel metal2 3818 7582 3818 7582 0 game.ballX\[5\]
rlabel metal1 2622 13974 2622 13974 0 game.ballX\[6\]
rlabel metal1 2714 14518 2714 14518 0 game.ballX\[7\]
rlabel metal2 6670 14654 6670 14654 0 game.ballX\[8\]
rlabel metal1 24564 7378 24564 7378 0 game.ballY\[0\]
rlabel metal2 23966 11424 23966 11424 0 game.ballY\[1\]
rlabel metal1 20102 8602 20102 8602 0 game.ballY\[2\]
rlabel metal1 20148 9146 20148 9146 0 game.ballY\[3\]
rlabel metal2 19550 10064 19550 10064 0 game.ballY\[4\]
rlabel metal1 17112 7922 17112 7922 0 game.ballY\[5\]
rlabel metal2 13846 6596 13846 6596 0 game.ballY\[6\]
rlabel metal2 13202 7548 13202 7548 0 game.ballY\[7\]
rlabel metal1 17516 19822 17516 19822 0 game.blue
rlabel metal1 10672 20298 10672 20298 0 game.col0
rlabel metal2 16514 18972 16514 18972 0 game.green
rlabel metal1 17894 19380 17894 19380 0 game.h\[0\]
rlabel metal1 15594 18734 15594 18734 0 game.h\[1\]
rlabel metal1 9568 12818 9568 12818 0 game.h\[2\]
rlabel metal1 8556 18258 8556 18258 0 game.h\[3\]
rlabel metal2 17618 17357 17618 17357 0 game.h\[4\]
rlabel metal1 7314 16660 7314 16660 0 game.h\[5\]
rlabel metal2 7038 17102 7038 17102 0 game.h\[6\]
rlabel metal1 5474 17272 5474 17272 0 game.h\[7\]
rlabel metal1 2530 14382 2530 14382 0 game.h\[8\]
rlabel metal1 10626 16524 10626 16524 0 game.h\[9\]
rlabel metal1 14582 12716 14582 12716 0 game.hit
rlabel metal1 4094 20026 4094 20026 0 game.hsync
rlabel metal1 8142 12920 8142 12920 0 game.inBallX
rlabel metal1 18262 12138 18262 12138 0 game.inBallY
rlabel metal2 18354 14144 18354 14144 0 game.inPaddle
rlabel metal1 15801 12818 15801 12818 0 game.new_game_n
rlabel metal1 10718 14994 10718 14994 0 game.offset\[0\]
rlabel metal1 18676 20434 18676 20434 0 game.offset\[1\]
rlabel metal2 19550 17986 19550 17986 0 game.offset\[2\]
rlabel metal1 13524 19346 13524 19346 0 game.offset\[3\]
rlabel metal1 11040 12818 11040 12818 0 game.offset\[4\]
rlabel metal2 28934 14654 28934 14654 0 game.paddle\[0\]
rlabel viali 26176 12818 26176 12818 0 game.paddle\[1\]
rlabel metal1 27784 7922 27784 7922 0 game.paddle\[2\]
rlabel via1 24994 10030 24994 10030 0 game.paddle\[3\]
rlabel metal2 28014 10846 28014 10846 0 game.paddle\[4\]
rlabel metal2 29210 10914 29210 10914 0 game.paddle\[5\]
rlabel metal1 29670 12682 29670 12682 0 game.paddle\[6\]
rlabel metal2 24334 13090 24334 13090 0 game.paddle\[7\]
rlabel metal1 23811 12818 23811 12818 0 game.paddle\[8\]
rlabel metal2 26542 14450 26542 14450 0 game.pause_n
rlabel metal1 15226 20332 15226 20332 0 game.red
rlabel metal1 13708 20434 13708 20434 0 game.row0
rlabel via3 13731 19380 13731 19380 0 game.speaker
rlabel metal1 31648 18734 31648 18734 0 game.up_key_n
rlabel metal2 14582 17255 14582 17255 0 game.v\[0\]
rlabel metal2 19274 17357 19274 17357 0 game.v\[1\]
rlabel metal1 28290 16116 28290 16116 0 game.v\[2\]
rlabel metal1 27094 17510 27094 17510 0 game.v\[3\]
rlabel metal1 24886 17034 24886 17034 0 game.v\[4\]
rlabel metal2 24794 16864 24794 16864 0 game.v\[5\]
rlabel metal2 15318 14110 15318 14110 0 game.v\[6\]
rlabel metal1 15226 13838 15226 13838 0 game.v\[7\]
rlabel metal1 20884 12682 20884 12682 0 game.v\[8\]
rlabel metal1 21482 14586 21482 14586 0 game.v\[9\]
rlabel metal2 17526 18394 17526 18394 0 game.vsync
rlabel metal1 12834 19414 12834 19414 0 lzc.a
rlabel metal2 31878 17034 31878 17034 0 net1
rlabel metal4 4508 21525 4508 21525 0 net10
rlabel metal4 3772 19757 3772 19757 0 net11
rlabel metal4 3036 21525 3036 21525 0 net12
rlabel via2 1794 19499 1794 19499 0 net13
rlabel metal4 1564 19757 1564 19757 0 net14
rlabel metal1 29608 19754 29608 19754 0 net15
rlabel metal1 30206 19414 30206 19414 0 net16
rlabel metal1 31341 17578 31341 17578 0 net17
rlabel metal1 30482 17238 30482 17238 0 net18
rlabel metal1 31924 19822 31924 19822 0 net2
rlabel metal1 26864 20026 26864 20026 0 net3
rlabel metal1 29762 18938 29762 18938 0 net4
rlabel metal2 28106 19380 28106 19380 0 net5
rlabel metal1 15502 20434 15502 20434 0 net6
rlabel metal1 4278 20332 4278 20332 0 net7
rlabel metal1 4048 20434 4048 20434 0 net8
rlabel metal1 3818 20502 3818 20502 0 net9
rlabel metal1 29056 20502 29056 20502 0 new_game.d
rlabel metal1 29164 20366 29164 20366 0 new_game.dff1
rlabel via1 30962 18666 30962 18666 0 pause.d
rlabel metal1 28658 18258 28658 18258 0 pause.dff1
rlabel metal2 18814 19516 18814 19516 0 qb
rlabel metal1 16238 19482 16238 19482 0 qg
rlabel metal1 16974 19346 16974 19346 0 qr
rlabel metal2 31878 19533 31878 19533 0 rst_n
rlabel metal4 30268 19281 30268 19281 0 ui_in[0]
rlabel metal4 29532 21525 29532 21525 0 ui_in[1]
rlabel metal4 28796 21525 28796 21525 0 ui_in[2]
rlabel metal4 28060 21525 28060 21525 0 ui_in[3]
rlabel metal4 27324 21321 27324 21321 0 ui_in[4]
rlabel metal4 12604 21389 12604 21389 0 uio_out[0]
rlabel metal4 11868 21457 11868 21457 0 uio_out[1]
rlabel metal2 13570 19210 13570 19210 0 uio_out[2]
rlabel metal1 11408 18870 11408 18870 0 uio_out[3]
rlabel metal1 8602 20502 8602 20502 0 uio_out[4]
rlabel metal2 9522 20723 9522 20723 0 uio_out[5]
rlabel metal1 13501 19958 13501 19958 0 uio_out[6]
rlabel via2 8142 20587 8142 20587 0 uio_out[7]
rlabel via2 18630 19499 18630 19499 0 uo_out[0]
rlabel via2 17066 20587 17066 20587 0 uo_out[1]
rlabel metal1 17112 19482 17112 19482 0 uo_out[2]
rlabel metal4 16284 21525 16284 21525 0 uo_out[3]
rlabel via2 16146 20587 16146 20587 0 uo_out[4]
rlabel metal1 13892 20026 13892 20026 0 uo_out[5]
rlabel metal4 14076 21525 14076 21525 0 uo_out[6]
rlabel via2 13570 20587 13570 20587 0 uo_out[7]
rlabel metal1 28708 19346 28708 19346 0 up_key.d
rlabel metal2 28382 19652 28382 19652 0 up_key.dff1
<< properties >>
string FIXED_BBOX 0 0 33580 21760
<< end >>
