`default_nettype none
`timescale 1ns/1ns
module hvsync_generator(
    input wire clk,
    input wire reset,
    output reg [9:0] sx,
    output reg [9:0] sy,
    output wire hsync,
    output wire vsync,
    output wire de
);
    // horizontal timings
    parameter HA_END = 639;           // end of active pixels
    parameter HS_STA = HA_END + 16;   // sync starts after front porch
    parameter HS_END = HS_STA + 96;   // sync ends
    parameter LINE   = 799;           // last pixel on line (after back porch)

    // vertical timings
    parameter VA_END = 479;           // end of active pixels
    parameter VS_STA = VA_END + 10;   // sync starts after front porch
    parameter VS_END = VS_STA + 2;    // sync ends
    parameter SCREEN = 524;           // last line on screen (after back porch)

    assign hsync = ~(sx >= HS_STA && sx < HS_END);
    assign vsync = ~(sy >= VS_STA && sy < VS_END);
    assign de = (sx <= HA_END && sy <= VA_END);

    always @(posedge clk) begin
        if (reset) begin
            sx <= 0;
            sy <= 0;
        end else begin
            if (sx == LINE) begin
                sx <= 0;
                sy <= (sy == SCREEN) ? 0 : sy + 1;
            end else begin
                sx <= sx + 1;
            end
        end
    end
endmodule
