magic
tech sky130A
magscale 1 2
timestamp 1713041211
<< nwell >>
rect -683 -419 683 419
<< pmos >>
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
<< pdiff >>
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
<< pdiffc >>
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
<< nsubdiff >>
rect -647 349 -551 383
rect 551 349 647 383
rect -647 287 -613 349
rect 613 287 647 349
rect -647 -349 -613 -287
rect 613 -349 647 -287
rect -647 -383 647 -349
<< nsubdiffcont >>
rect -551 349 551 383
rect -647 -287 -613 287
rect 613 -287 647 287
<< poly >>
rect -487 281 -287 297
rect -487 247 -471 281
rect -303 247 -287 281
rect -487 200 -287 247
rect -229 281 -29 297
rect -229 247 -213 281
rect -45 247 -29 281
rect -229 200 -29 247
rect 29 281 229 297
rect 29 247 45 281
rect 213 247 229 281
rect 29 200 229 247
rect 287 281 487 297
rect 287 247 303 281
rect 471 247 487 281
rect 287 200 487 247
rect -487 -247 -287 -200
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -487 -297 -287 -281
rect -229 -247 -29 -200
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect -229 -297 -29 -281
rect 29 -247 229 -200
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 29 -297 229 -281
rect 287 -247 487 -200
rect 287 -281 303 -247
rect 471 -281 487 -247
rect 287 -297 487 -281
<< polycont >>
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
<< locali >>
rect -647 349 -551 383
rect 551 349 647 383
rect 613 287 647 349
rect -303 247 -287 281
rect -45 247 -29 281
rect 213 247 229 281
rect 471 247 487 281
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect -303 -281 -287 -247
rect -45 -281 -29 -247
rect 213 -281 229 -247
rect 471 -281 487 -247
rect 613 -349 647 -287
rect -647 -383 647 -349
<< viali >>
rect -647 287 -613 349
rect -647 -287 -613 287
rect -488 247 -471 281
rect -471 247 -320 281
rect -230 247 -213 281
rect -213 247 -62 281
rect 28 247 45 281
rect 45 247 196 281
rect 286 247 303 281
rect 303 247 454 281
rect -533 21 -499 171
rect -275 -171 -241 -21
rect -17 21 17 171
rect 241 -171 275 -21
rect 499 21 533 171
rect -488 -281 -471 -247
rect -471 -281 -320 -247
rect -230 -281 -213 -247
rect -213 -281 -62 -247
rect 28 -281 45 -247
rect 45 -281 196 -247
rect 286 -281 303 -247
rect 303 -281 454 -247
rect -647 -349 -613 -287
<< metal1 >>
rect -653 349 -607 361
rect -653 -349 -647 349
rect -613 -349 -607 349
rect -500 281 -308 287
rect -500 247 -488 281
rect -320 247 -308 281
rect -500 241 -308 247
rect -242 281 -50 287
rect -242 247 -230 281
rect -62 247 -50 281
rect -242 241 -50 247
rect 16 281 208 287
rect 16 247 28 281
rect 196 247 208 281
rect 16 241 208 247
rect 274 281 466 287
rect 274 247 286 281
rect 454 247 466 281
rect 274 241 466 247
rect -539 171 -493 183
rect -539 21 -533 171
rect -499 21 -493 171
rect -539 9 -493 21
rect -23 171 23 183
rect -23 21 -17 171
rect 17 21 23 171
rect -23 9 23 21
rect 493 171 539 183
rect 493 21 499 171
rect 533 21 539 171
rect 493 9 539 21
rect -281 -21 -235 -9
rect -281 -171 -275 -21
rect -241 -171 -235 -21
rect -281 -183 -235 -171
rect 235 -21 281 -9
rect 235 -171 241 -21
rect 275 -171 281 -21
rect 235 -183 281 -171
rect -500 -247 -308 -241
rect -500 -281 -488 -247
rect -320 -281 -308 -247
rect -500 -287 -308 -281
rect -242 -247 -50 -241
rect -242 -281 -230 -247
rect -62 -281 -50 -247
rect -242 -287 -50 -281
rect 16 -247 208 -241
rect 16 -281 28 -247
rect 196 -281 208 -247
rect 16 -287 208 -281
rect 274 -247 466 -241
rect 274 -281 286 -247
rect 454 -281 466 -247
rect 274 -287 466 -281
rect -653 -361 -607 -349
<< properties >>
string FIXED_BBOX -630 -366 630 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate -100 viagb 0 viagr 0 viagl 100 viagt 0
<< end >>
