magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -1199 -410 1199 410
<< nmos >>
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
<< ndiff >>
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
<< ndiffc >>
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
<< psubdiff >>
rect -1163 340 -1067 374
rect 1067 340 1163 374
rect -1163 278 -1129 340
rect 1129 278 1163 340
rect -1163 -340 -1129 -278
rect 1129 -340 1163 -278
rect -1163 -374 1163 -340
<< psubdiffcont >>
rect -1067 340 1067 374
rect -1163 -278 -1129 278
rect 1129 -278 1163 278
<< poly >>
rect -1003 272 -803 288
rect -1003 238 -987 272
rect -819 238 -803 272
rect -1003 200 -803 238
rect -745 272 -545 288
rect -745 238 -729 272
rect -561 238 -545 272
rect -745 200 -545 238
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect 545 272 745 288
rect 545 238 561 272
rect 729 238 745 272
rect 545 200 745 238
rect 803 272 1003 288
rect 803 238 819 272
rect 987 238 1003 272
rect 803 200 1003 238
rect -1003 -238 -803 -200
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -1003 -288 -803 -272
rect -745 -238 -545 -200
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -745 -288 -545 -272
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
rect 545 -238 745 -200
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 545 -288 745 -272
rect 803 -238 1003 -200
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect 803 -288 1003 -272
<< polycont >>
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
<< locali >>
rect -1163 278 -1129 374
rect 1129 278 1163 374
rect -1003 238 -987 272
rect -819 238 -803 272
rect -745 238 -729 272
rect -561 238 -545 272
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect 545 238 561 272
rect 729 238 745 272
rect 803 238 819 272
rect 987 238 1003 272
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect -1163 -374 1163 -340
<< viali >>
rect -1129 340 -1067 374
rect -1067 340 1067 374
rect 1067 340 1129 374
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect -1163 -278 -1129 -68
rect -1049 21 -1015 171
rect -791 -171 -757 -21
rect -533 21 -499 171
rect -275 -171 -241 -21
rect -17 21 17 171
rect 241 -171 275 -21
rect 499 21 533 171
rect 757 -171 791 -21
rect 1015 21 1049 171
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
rect -1163 -340 -1129 -278
rect 1129 -278 1163 -68
rect 1129 -340 1163 -278
<< metal1 >>
rect -1141 374 1141 380
rect -1141 340 -1129 374
rect 1129 340 1141 374
rect -1141 334 1141 340
rect -999 272 -807 278
rect -999 238 -987 272
rect -819 238 -807 272
rect -999 232 -807 238
rect -741 272 -549 278
rect -741 238 -729 272
rect -561 238 -549 272
rect -741 232 -549 238
rect -483 272 -291 278
rect -483 238 -471 272
rect -303 238 -291 272
rect -483 232 -291 238
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect 291 272 483 278
rect 291 238 303 272
rect 471 238 483 272
rect 291 232 483 238
rect 549 272 741 278
rect 549 238 561 272
rect 729 238 741 272
rect 549 232 741 238
rect 807 272 999 278
rect 807 238 819 272
rect 987 238 999 272
rect 807 232 999 238
rect -1055 171 -1009 183
rect -1055 21 -1049 171
rect -1015 21 -1009 171
rect -1055 9 -1009 21
rect -539 171 -493 183
rect -539 21 -533 171
rect -499 21 -493 171
rect -539 9 -493 21
rect -23 171 23 183
rect -23 21 -17 171
rect 17 21 23 171
rect -23 9 23 21
rect 493 171 539 183
rect 493 21 499 171
rect 533 21 539 171
rect 493 9 539 21
rect 1009 171 1055 183
rect 1009 21 1015 171
rect 1049 21 1055 171
rect 1009 9 1055 21
rect -797 -21 -751 -9
rect -1169 -68 -1123 -56
rect -1169 -340 -1163 -68
rect -1129 -340 -1123 -68
rect -797 -171 -791 -21
rect -757 -171 -751 -21
rect -797 -183 -751 -171
rect -281 -21 -235 -9
rect -281 -171 -275 -21
rect -241 -171 -235 -21
rect -281 -183 -235 -171
rect 235 -21 281 -9
rect 235 -171 241 -21
rect 275 -171 281 -21
rect 235 -183 281 -171
rect 751 -21 797 -9
rect 751 -171 757 -21
rect 791 -171 797 -21
rect 751 -183 797 -171
rect 1123 -68 1169 -56
rect -999 -238 -807 -232
rect -999 -272 -987 -238
rect -819 -272 -807 -238
rect -999 -278 -807 -272
rect -741 -238 -549 -232
rect -741 -272 -729 -238
rect -561 -272 -549 -238
rect -741 -278 -549 -272
rect -483 -238 -291 -232
rect -483 -272 -471 -238
rect -303 -272 -291 -238
rect -483 -278 -291 -272
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
rect 291 -238 483 -232
rect 291 -272 303 -238
rect 471 -272 483 -238
rect 291 -278 483 -272
rect 549 -238 741 -232
rect 549 -272 561 -238
rect 729 -272 741 -238
rect 549 -278 741 -272
rect 807 -238 999 -232
rect 807 -272 819 -238
rect 987 -272 999 -238
rect 807 -278 999 -272
rect -1169 -352 -1123 -340
rect 1123 -340 1129 -68
rect 1163 -340 1169 -68
rect 1123 -352 1169 -340
<< properties >>
string FIXED_BBOX -1146 -357 1146 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
