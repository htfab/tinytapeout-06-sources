magic
tech sky130A
magscale 1 2
timestamp 1713420874
<< locali >>
rect 1052 2536 3482 2578
rect 1052 2370 1396 2536
rect 3258 2370 3482 2536
rect 1052 2290 3482 2370
rect 1056 534 2110 2196
rect 2404 534 3478 2184
rect 1056 196 3478 534
rect 1056 184 2110 196
rect 1056 -330 1206 184
rect 3242 -330 3478 196
rect 1056 -416 3478 -330
rect 1052 -468 3478 -416
rect 1052 -702 1230 -468
rect 1048 -852 1230 -702
rect 3292 -852 3478 -468
rect 1048 -958 3478 -852
<< viali >>
rect 1396 2370 3258 2536
rect 1230 -852 3292 -468
<< metal1 >>
rect 1120 2536 3360 2572
rect 1120 2370 1396 2536
rect 3258 2370 3360 2536
rect 1120 2338 3360 2370
rect 2174 1622 2376 2338
rect 2166 916 2354 1134
rect 2166 570 3478 916
rect 2166 364 2354 570
rect 1654 254 2804 364
rect 1648 252 2804 254
rect 1648 184 2812 252
rect 1504 88 1544 96
rect 1648 88 1900 184
rect 1962 88 2002 108
rect 1192 -156 1202 44
rect 1402 -156 1412 44
rect 1504 40 2002 88
rect 1504 -160 1660 40
rect 1860 -160 2002 40
rect 2424 96 2464 108
rect 2560 96 2812 184
rect 2888 96 2928 108
rect 2424 40 2928 96
rect 1504 -206 2002 -160
rect 2108 -164 2118 36
rect 2318 -164 2328 36
rect 2424 -160 2570 40
rect 2770 -160 2928 40
rect 3018 -160 3028 40
rect 3228 -160 3238 40
rect 2424 -206 2928 -160
rect 1504 -218 1974 -206
rect 2446 -214 2896 -206
rect 1524 -222 1974 -218
rect 1154 -468 3384 -374
rect 1154 -852 1230 -468
rect 3292 -852 3384 -468
rect 1154 -922 3384 -852
<< via1 >>
rect 1202 -156 1402 44
rect 1660 -160 1860 40
rect 2118 -164 2318 36
rect 2570 -160 2770 40
rect 3028 -160 3228 40
rect 1296 -498 3148 -478
rect 1280 -644 3152 -498
<< metal2 >>
rect 1202 44 1402 54
rect 1202 -166 1402 -156
rect 1660 40 1860 50
rect 1252 -438 1360 -166
rect 1660 -170 1860 -160
rect 2118 36 2318 46
rect 2118 -174 2318 -164
rect 2570 40 2770 50
rect 2570 -170 2770 -160
rect 3028 40 3228 50
rect 3028 -170 3228 -160
rect 2164 -438 2272 -174
rect 3074 -438 3182 -170
rect 1246 -478 3210 -438
rect 1246 -498 1296 -478
rect 3148 -498 3210 -478
rect 1246 -644 1280 -498
rect 3152 -644 3210 -498
rect 1246 -686 3210 -644
use sky130_fd_pr__nfet_01v8_VWWVRL  XM6
timestamp 1713420874
transform 1 0 2221 0 1 -60
box -1083 -310 1083 310
use sky130_fd_pr__res_xhigh_po_0p35_5BGKUX  XR1
timestamp 1713420874
transform 1 0 2261 0 1 1356
box -201 -862 201 862
<< labels >>
flabel metal1 2146 2360 2346 2560 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 2184 -922 2384 -722 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 3238 654 3438 854 0 FreeSans 256 0 0 0 VBIAS
port 2 nsew
<< end >>
