* NGSPICE file created from tt_um_argunda_tiny_opamp.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_5BGKUX a_n35_n696# a_n165_n826# a_n35_264#
X0 a_n35_264# a_n35_n696# a_n165_n826# sky130_fd_pr__res_xhigh_po_0p35 l=2.8
.ends

.subckt sky130_fd_pr__nfet_01v8_VWWVRL a_n29_n100# a_887_n100# a_429_n100# a_n887_n188#
+ a_n1047_n274# a_n429_n188# a_487_n188# a_n945_n100# a_29_n188# a_n487_n100#
X0 a_887_n100# a_487_n188# a_429_n100# a_n1047_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=11600,516
X1 a_429_n100# a_29_n188# a_n29_n100# a_n1047_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X2 a_n487_n100# a_n887_n188# a_n945_n100# a_n1047_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=5800,258
X3 a_n29_n100# a_n429_n188# a_n487_n100# a_n1047_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
.ends

.subckt vbias_resistor VDD VBIAS VSS
XXR1 VBIAS VSS VDD sky130_fd_pr__res_xhigh_po_0p35_5BGKUX
XXM6 VSS VSS VBIAS VBIAS VSS VBIAS VBIAS VSS VBIAS VBIAS sky130_fd_pr__nfet_01v8_VWWVRL
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_8TELWR a_n108_n250# a_n50_n338# a_n210_n424# a_50_n250#
X0 a_50_n250# a_n50_n338# a_n108_n250# a_n210_n424# sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
**devattr s=29000,1116 d=29000,1116
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GW6ZVV a_n887_n197# a_1345_n100# a_n29_n100# a_945_n197#
+ a_887_n100# a_n429_n197# a_487_n197# a_429_n100# a_29_n197# a_n1403_n100# w_n1541_n319#
+ a_n1345_n197# a_n945_n100# a_n487_n100#
X0 a_1345_n100# a_945_n197# a_887_n100# w_n1541_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=11600,516
X1 a_429_n100# a_29_n197# a_n29_n100# w_n1541_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X2 a_n487_n100# a_n887_n197# a_n945_n100# w_n1541_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X3 a_n29_n100# a_n429_n197# a_n487_n100# w_n1541_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X4 a_n945_n100# a_n1345_n197# a_n1403_n100# w_n1541_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=5800,258
X5 a_887_n100# a_487_n197# a_429_n100# w_n1541_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
.ends

.subckt sky130_fd_pr__nfet_01v8_WWWVRA a_n258_n100# a_1574_n100# a_1116_n100# a_n200_n188#
+ a_658_n100# a_n1574_n188# a_n1116_n188# a_n1734_n274# a_n1632_n100# a_1174_n188#
+ a_n658_n188# a_n1174_n100# a_716_n188# a_258_n188# a_200_n100# a_n716_n100#
X0 a_200_n100# a_n200_n188# a_n258_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X1 a_n1174_n100# a_n1574_n188# a_n1632_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=5800,258
X2 a_n258_n100# a_n658_n188# a_n716_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X3 a_n716_n100# a_n1116_n188# a_n1174_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X4 a_658_n100# a_258_n188# a_200_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X5 a_1574_n100# a_1174_n188# a_1116_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=11600,516
X6 a_1116_n100# a_716_n188# a_658_n100# a_n1734_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_ER3WAW a_1293_n197# a_n761_n197# a_1235_n100#
+ a_n1551_n197# a_761_n100# a_n29_n100# a_1393_n100# a_1451_n197# a_n187_n100# a_1551_n100#
+ a_n819_n100# a_n345_n100# a_n1609_n100# a_29_n197# a_n977_n100# a_n1135_n100# a_n129_n197#
+ a_187_n197# w_n1747_n319# a_129_n100# a_n503_n100# a_n1293_n100# a_n287_n197# a_819_n197#
+ a_n661_n100# a_345_n197# a_n1077_n197# a_287_n100# a_n1451_n100# a_n919_n197# a_977_n197#
+ a_n445_n197# a_919_n100# a_503_n197# a_n1235_n197# a_445_n100# a_1077_n100# a_1135_n197#
+ a_n603_n197# a_n1393_n197# a_661_n197# a_603_n100#
X0 a_n1293_n100# a_n1393_n197# a_n1451_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X1 a_n1451_n100# a_n1551_n197# a_n1609_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
**devattr s=11600,516 d=5800,258
X2 a_n977_n100# a_n1077_n197# a_n1135_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X3 a_n1135_n100# a_n1235_n197# a_n1293_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X4 a_n661_n100# a_n761_n197# a_n819_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X5 a_129_n100# a_29_n197# a_n29_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X6 a_n187_n100# a_n287_n197# a_n345_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X7 a_n819_n100# a_n919_n197# a_n977_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X8 a_n345_n100# a_n445_n197# a_n503_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X9 a_n503_n100# a_n603_n197# a_n661_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X10 a_n29_n100# a_n129_n197# a_n187_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X11 a_1393_n100# a_1293_n197# a_1235_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X12 a_1077_n100# a_977_n197# a_919_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X13 a_1551_n100# a_1451_n197# a_1393_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=11600,516
X14 a_761_n100# a_661_n197# a_603_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X15 a_287_n100# a_187_n197# a_129_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X16 a_1235_n100# a_1135_n197# a_1077_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X17 a_445_n100# a_345_n197# a_287_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X18 a_919_n100# a_819_n197# a_761_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X19 a_603_n100# a_503_n197# a_445_n100# w_n1747_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
.ends

.subckt opamp VBIAS VDD MINUS PLUS VOUT VSS
XXM1 V1 PLUS VSS m1_2578_n2492# sky130_fd_pr__nfet_01v8_lvt_8TELWR
XXM2 V2 MINUS VSS m1_2578_n2492# sky130_fd_pr__nfet_01v8_lvt_8TELWR
XXM3 VSS VSS m1_2578_n2492# VBIAS VSS VBIAS VBIAS VSS VBIAS m1_2578_n2492# sky130_fd_pr__nfet_01v8_VWWVRL
XXM4 V2 VDD V2 V2 V2 V2 V2 VDD V2 VDD VDD V2 V2 VDD sky130_fd_pr__pfet_01v8_lvt_GW6ZVV
XXM5 V2 VDD V1 V2 V1 V2 V2 VDD V2 VDD VDD V2 V1 VDD sky130_fd_pr__pfet_01v8_lvt_GW6ZVV
XXM7 VSS VSS VOUT VBIAS VSS VBIAS VBIAS VSS VOUT VBIAS VBIAS VSS VBIAS VBIAS VOUT
+ VOUT sky130_fd_pr__nfet_01v8_WWWVRA
XXM8 V1 V1 VOUT V1 VDD VOUT VDD V1 VDD VOUT VDD VOUT VOUT V1 VOUT VDD V1 V1 VDD VDD
+ VDD VOUT V1 V1 VOUT V1 V1 VOUT VDD V1 V1 V1 VOUT V1 V1 VDD VDD V1 V1 V1 V1 VOUT
+ sky130_fd_pr__pfet_01v8_lvt_ER3WAW
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=4.73
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=4.73
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=2.89
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=2.89
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=1.05
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.05
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12054 ps=1.304827 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12353 pd=1.162647 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.193015 ps=1.816635 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.081066 ps=0.762987 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193015 pd=1.816635 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.081066 pd=0.762987 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0.118685 ps=1.284752 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.144761 ps=1.362476 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.077887 ps=0.843119 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.081066 pd=0.762987 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12353 ps=1.162647 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.12054 pd=1.304827 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0.077887 ps=0.843119 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=1.97
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.97
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.943333 as=0.1525 ps=1.305 w=1 l=0.15
**devattr s=6100,261 d=10400,504
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4030,192
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=4030,192 d=3510,184
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.943333 as=0.28 ps=2.56 w=1 l=0.15
**devattr s=11200,512 d=13100,331
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.305 ps=1.943333 w=1 l=0.15
**devattr s=13100,331 d=7800,278
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=6100,261
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073937 pd=0.752655 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073937 pd=0.752655 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103351 pd=0.894953 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.073937 ps=0.752655 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.17604 ps=1.792035 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.159949 ps=1.385047 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VPB VNB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2940,154
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.088214 pd=0.825097 as=0.082425 ps=0.8125 w=0.42 l=0.15
**devattr s=2646,147 d=5630,265
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.137852 ps=1.465772 w=0.65 l=0.15
**devattr s=4136,200 d=6760,364
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.088214 pd=0.825097 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.089074 pd=0.947114 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=4136,200
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.210032 ps=1.964516 w=1 l=0.15
**devattr s=5630,265 d=10400,504
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.088214 pd=0.825097 as=0.082425 ps=0.8125 w=0.42 l=0.15
**devattr s=3948,178 d=5124,206
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.082425 pd=0.8125 as=0.088214 ps=0.825097 w=0.42 l=0.15
**devattr s=5124,206 d=2646,147
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.082425 pd=0.8125 as=0.088214 ps=0.825097 w=0.42 l=0.15
**devattr s=2268,138 d=3948,178
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
**devattr s=2940,154 d=2436,142
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.089074 pd=0.947114 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.102877 pd=0.95413 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.244946 ps=2.271739 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.087768 pd=0.816449 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.102877 ps=0.95413 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.135832 ps=1.263551 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=0.59
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=0.59
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.187633 pd=1.713333 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=6400,264 d=6200,262
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
**devattr s=2990,176 d=6760,364
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.11375 ps=1 w=0.65 l=0.15
**devattr s=4550,200 d=4030,192
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.187633 ps=1.713333 w=1 l=0.15
**devattr s=6200,262 d=10400,504
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.256425 pd=2.52 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=5400,254 d=10114,504
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.187633 ps=1.713333 w=1 l=0.15
**devattr s=10116,504 d=6400,264
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4550,200
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=4030,192 d=6760,364
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.256425 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=6760,364 d=2990,176
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111244 pd=0.929204 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.264867 ps=2.212389 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13602 ps=1.457047 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.111244 ps=0.929204 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111244 pd=0.929204 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08789 pd=0.941476 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08789 ps=0.941476 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213258 pd=1.962121 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10600,506
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.213258 ps=1.962121 w=1 l=0.15
**devattr s=5960,265 d=5400,254
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.136485 pd=1.255758 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=5960,265
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138408 ps=1.428488 w=0.65 l=0.15
**devattr s=3880,195 d=3510,184
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.138408 pd=1.428488 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.089433 pd=0.923023 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3475 ps=2.195 w=1 l=0.15
**devattr s=14600,346 d=4200,242
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3475 ps=2.195 w=1 l=0.15
**devattr s=12000,520 d=5400,254
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=2730,172
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=7800,380
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=3510,184
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3475 pd=2.195 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=14600,346
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3475 pd=2.195 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=14400,544
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6600,266
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.127256 ps=1.376226 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.203665 pd=1.928458 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.130345 pd=1.234213 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.203665 ps=1.928458 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.085539 ps=0.809952 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.082227 pd=0.889254 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.127256 pd=1.376226 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.203665 pd=1.928458 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.085539 pd=0.809952 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0.125298 ps=1.355053 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.152748 ps=1.446343 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.082227 pd=0.889254 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.082227 ps=0.889254 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.085539 pd=0.809952 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.130345 ps=1.234213 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.127256 pd=1.376226 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0.082227 ps=0.889254 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.082227 pd=0.889254 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.084613 pd=0.797257 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.084613 ps=0.797257 w=0.42 l=0.15
**devattr s=2772,150 d=4704,280
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.084613 ps=0.797257 w=0.42 l=0.15
**devattr s=6334,279 d=3066,157
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.113356 pd=0.947749 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5796,222
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7728,268
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.113356 ps=0.947749 w=0.42 l=0.15
**devattr s=5796,222 d=4368,272
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=1764,126
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113356 ps=0.947749 w=0.42 l=0.15
**devattr s=4514,209 d=2772,150
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20146 pd=1.89823 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=6334,279
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.175432 pd=1.466754 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4514,209
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
.ends

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.087298 pd=0.938658 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.087298 ps=0.938658 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135104 ps=1.452685 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.086218 pd=0.789718 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.205282 ps=1.880282 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VPB VNB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.139399 ps=0.987313 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.331903 ps=2.350746 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.139399 ps=0.987313 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139399 pd=0.987313 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.154085 pd=1.044112 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139399 pd=0.987313 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.238465 ps=1.615888 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=3835,189
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=5900,259 d=10600,506
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=3640,186
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=5900,259
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
**devattr s=3835,189 d=6890,366
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.163583 pd=1.37 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=6760,364
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.544 as=0.172 ps=1.544 w=1 l=0.15
**devattr s=6600,266 d=6600,266
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.544 as=0.172 ps=1.544 w=1 l=0.15
**devattr s=5400,254 d=6600,266
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.544 as=0.172 ps=1.544 w=1 l=0.15
**devattr s=6600,266 d=10400,504
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.544 as=0.172 ps=1.544 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
**devattr s=7345,243 d=3510,184
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.544 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.544 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.163583 ps=1.37 w=0.65 l=0.15
**devattr s=6435,229 d=7345,243
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.163583 pd=1.37 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6435,229
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
.ends

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.141375 ps=1.41 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.003333 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
**devattr s=9400,294 d=4200,242
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.003333 as=0.28 ps=2.56 w=1 l=0.15
**devattr s=11200,512 d=14900,349
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.141375 ps=1.41 w=0.65 l=0.15
**devattr s=4550,200 d=3510,184
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
**devattr s=4700,247 d=9400,294
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.41 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.41 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=4550,200
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.335 ps=2.003333 w=1 l=0.15
**devattr s=14900,349 d=4700,247
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.3375 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6900,269
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.16875 ps=1.3375 w=1 l=0.15
**devattr s=6900,269 d=6400,264
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4290,196
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.144083 ps=1.31 w=0.65 l=0.15
**devattr s=4485,199 d=4160,194
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.144083 pd=1.31 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=4485,199
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.144083 pd=1.31 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=8320,388
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.3375 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6600,266
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=12800,528
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.16875 ps=1.3375 w=1 l=0.15
**devattr s=6600,266 d=6600,266
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.118083 ps=1.23 w=0.65 l=0.15
**devattr s=3640,186 d=5070,208
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.118083 ps=1.23 w=0.65 l=0.15
**devattr s=3640,186 d=3640,186
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.925 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.925 as=0.1575 ps=1.315 w=1 l=0.15
**devattr s=7000,270 d=6400,264
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.108875 ps=0.985 w=0.65 l=0.15
**devattr s=3640,186 d=3640,186
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1575 ps=1.315 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.118083 ps=1.23 w=0.65 l=0.15
**devattr s=6890,366 d=3640,186
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.2125 ps=1.925 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=7000,270
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2125 ps=1.925 w=1 l=0.15
**devattr s=6400,264 d=5600,256
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.108875 ps=0.985 w=0.65 l=0.15
**devattr s=5070,208 d=3640,186
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073388 pd=0.748938 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.067596 pd=0.732251 as=0.1092 ps=1.36 w=0.42 l=0.5
**devattr s=4368,272 d=3880,195
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.174735 ps=1.783186 w=1 l=0.15
**devattr s=5630,265 d=10400,504
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.067596 pd=0.732251 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073388 pd=0.748938 as=0.1092 ps=1.36 w=0.42 l=0.5
**devattr s=4368,272 d=5630,265
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.067596 ps=0.732251 w=0.42 l=0.5
**devattr s=2268,138 d=4368,272
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.073388 ps=0.748938 w=0.42 l=0.5
**devattr s=2268,138 d=4368,272
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.104613 ps=1.133246 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.204706 pd=1.635294 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6960,278
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.828235 as=0.143294 ps=1.144706 w=0.7 l=0.15
**devattr s=6960,278 d=7280,384
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.611765 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
.ends

.subckt sky130_fd_sc_hd__nand4_1 VPB VNB VPWR VGND A C D Y B
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.2075 ps=1.915 w=1 l=0.15
**devattr s=5400,254 d=6600,266
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.915 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6600,266 d=12000,520
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.915 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=7800,380
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.2075 ps=1.915 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.228583 ps=1.57 w=0.65 l=0.15
**devattr s=10270,288 d=3575,185
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5500,255
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.18 ps=1.693333 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.228583 pd=1.57 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=10270,288
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.228583 pd=1.57 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.18 ps=1.693333 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
**devattr s=3575,185 d=3640,186
.ends

.subckt sky130_fd_sc_hd__o211a_1 VNB VPB VGND VPWR X A1 A2 B1 C1
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.256667 as=0.151667 ps=1.333333 w=0.65 l=0.15
**devattr s=6760,364 d=4225,195
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.151667 ps=1.333333 w=0.65 l=0.15
**devattr s=5720,218 d=4550,200
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.246667 pd=1.826667 as=0.2175 ps=1.935 w=1 l=0.15
**devattr s=7000,270 d=12000,520
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.935 as=0.246667 ps=1.826667 w=1 l=0.15
**devattr s=8800,288 d=7000,270
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.246667 pd=1.826667 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6500,265 d=8800,288
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.2175 ps=1.935 w=1 l=0.15
**devattr s=10400,504 d=6500,265
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
**devattr s=4550,200 d=7800,380
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.935 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.256667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.151667 pd=1.333333 as=0.12675 ps=1.256667 w=0.65 l=0.15
**devattr s=4225,195 d=5720,218
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.208803 ps=1.887324 w=1 l=0.15
**devattr s=5930,268 d=11200,512
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.107931 ps=1.143456 w=0.65 l=0.15
**devattr s=4075,198 d=7280,372
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.087697 pd=0.792676 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.06974 ps=0.738848 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.06974 pd=0.738848 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.06974 pd=0.738848 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VNB VPB VGND VPWR X A2 A1 B1_N
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=5400,254
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.216269 ps=1.395992 w=0.65 l=0.15
**devattr s=5436,220 d=3510,184
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.189825 ps=1.883041 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.216269 ps=1.395992 w=0.65 l=0.15
**devattr s=10335,289 d=6760,364
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.079726 pd=0.790877 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.189825 ps=1.883041 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3640,186
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.139743 pd=0.902025 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=5436,220
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.189825 pd=1.883041 as=0.178333 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=5600,256
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.216269 pd=1.395992 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=10335,289
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.099715 ps=0.992215 w=0.42 l=0.15
**devattr s=4368,272 d=4314,272
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.189198 ps=2.018657 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.079463 ps=0.847836 w=0.42 l=0.15
**devattr s=4368,272 d=4348,272
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
**devattr s=4313,272 d=1764,126
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.079463 pd=0.847836 as=0.08575 ps=0.996667 w=0.42 l=0.15
**devattr s=2975,163 d=5689,267
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2142,135
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.15432 ps=1.53557 w=0.65 l=0.15
**devattr s=4891,216 d=6760,364
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08575 pd=0.996667 as=0.079463 ps=0.847836 w=0.42 l=0.15
**devattr s=2268,138 d=2975,163
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.079463 pd=0.847836 as=0.08575 ps=0.996667 w=0.42 l=0.15
**devattr s=4340,272 d=2268,138
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.099715 pd=0.992215 as=0.05355 ps=0.675 w=0.42 l=0.15
**devattr s=2142,135 d=4891,216
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.220489 ps=2.195652 w=1 l=0.15
**devattr s=5930,268 d=11000,510
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.081793 ps=0.928582 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.060375 pd=0.7075 as=0.081793 ps=0.928582 w=0.42 l=0.15
**devattr s=4368,272 d=2562,145
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.126585 ps=1.437091 w=0.65 l=0.15
**devattr s=4075,198 d=7150,370
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=1806,127
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
**devattr s=1806,127 d=2562,145
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.060375 pd=0.7075 as=0.081793 ps=0.928582 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092605 pd=0.922174 as=0.06405 ps=0.725 w=0.42 l=0.15
**devattr s=2562,145 d=5930,268
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2730,149
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.092605 ps=0.922174 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.081793 pd=0.928582 as=0.060375 ps=0.7075 w=0.42 l=0.15
**devattr s=2562,145 d=2268,138
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.081793 pd=0.928582 as=0.060375 ps=0.7075 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VNB VPB VGND VPWR B1_N A1 A2 X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066633 ps=0.67519 w=0.42 l=0.15
**devattr s=4010,197 d=4368,272
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.278216 pd=2.336257 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=11200,512
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.103122 pd=1.044937 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4010,197
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.116851 ps=0.981228 w=0.42 l=0.15
**devattr s=7430,283 d=4704,280
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103122 pd=1.044937 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.278216 ps=2.336257 w=1 l=0.15
**devattr s=12000,520 d=6600,266
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.103122 ps=1.044937 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.278216 pd=2.336257 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=7430,283
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VPB VGND VPWR VNB B1 X D1 A1 A2 C1
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19435 pd=1.378 as=0.082875 ps=0.905 w=0.65 l=0.15
**devattr s=3315,181 d=7540,376
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.19435 pd=1.378 as=0.143 ps=1.09 w=0.65 l=0.15
**devattr s=4030,192 d=4680,202
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
**devattr s=5000,250 d=7200,272
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.19435 pd=1.378 as=0.2145 ps=1.96 w=0.65 l=0.15
**devattr s=8580,392 d=10985,299
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
**devattr s=15400,554 d=5000,250
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.283333 pd=1.9 as=0.18 ps=1.36 w=1 l=0.15
**devattr s=7200,272 d=11200,312
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.283333 pd=1.9 as=0.178333 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=11600,516
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.143 ps=1.09 w=0.65 l=0.15
**devattr s=7410,244 d=3315,181
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.19435 ps=1.378 w=0.65 l=0.15
**devattr s=10985,299 d=4030,192
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.283333 ps=1.9 w=1 l=0.15
**devattr s=11200,312 d=5400,254
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.19435 ps=1.378 w=0.65 l=0.15
**devattr s=4680,202 d=7410,244
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=10600,506
.ends

.subckt sky130_fd_sc_hd__and4_2 VNB VPB VGND VPWR X D C B A
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.206073 pd=1.674128 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=7800,380
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133155 pd=1.081744 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7006,253
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.305571 ps=2.383152 w=1 l=0.15
**devattr s=11198,323 d=6600,266
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
**devattr s=2478,143 d=3192,160
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.066675 pd=0.7375 as=0.12834 ps=1.000924 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305571 pd=2.383152 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=12000,520
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.066675 pd=0.7375 as=0.12834 ps=1.000924 w=0.42 l=0.15
**devattr s=4368,272 d=2982,155
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12834 pd=1.000924 as=0.066675 ps=0.7375 w=0.42 l=0.15
**devattr s=2352,140 d=11198,323
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.206073 ps=1.674128 w=0.65 l=0.15
**devattr s=7006,253 d=4290,196
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12834 pd=1.000924 as=0.066675 ps=0.7375 w=0.42 l=0.15
**devattr s=2982,155 d=3108,158
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2478,143
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2025 ps=1.905 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.131625 ps=1.38 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2025 pd=1.905 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.131625 pd=1.38 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.131625 ps=1.38 w=0.65 l=0.15
**devattr s=7280,372 d=3510,184
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.131625 pd=1.38 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2025 ps=1.905 w=1 l=0.15
**devattr s=11200,512 d=5400,254
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2025 pd=1.905 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138125 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.4 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.4 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138125 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
.ends

.subckt sky130_fd_sc_hd__a31oi_2 VNB VPB VPWR VGND B1 Y A1 A2 A3
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.143 ps=1.415 w=0.65 l=0.15
**devattr s=4680,202 d=4550,200
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226667 pd=1.453333 as=0.1775 ps=1.605 w=1 l=0.15
**devattr s=5400,254 d=16400,364
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.605 as=0.226667 ps=1.453333 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.605 as=0.175 ps=1.35 w=1 l=0.15
**devattr s=7000,270 d=10400,504
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.143 ps=1.415 w=0.65 l=0.15
**devattr s=6760,364 d=3900,190
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226667 pd=1.453333 as=0.1775 ps=1.605 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.605 as=0.226667 ps=1.453333 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.10075 ps=0.96 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.092625 ps=0.935 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.605 as=0.226667 ps=1.453333 w=1 l=0.15
**devattr s=16400,364 d=7200,272
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.1775 ps=1.605 w=1 l=0.15
**devattr s=7200,272 d=7000,270
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.415 as=0.10075 ps=0.96 w=0.65 l=0.15
**devattr s=4550,200 d=6760,364
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.415 as=0.092625 ps=0.935 w=0.65 l=0.15
**devattr s=3900,190 d=4680,202
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226667 pd=1.453333 as=0.1775 ps=1.605 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.076267 ps=0.849013 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.076267 ps=0.849013 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.076267 pd=0.849013 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.076267 pd=0.849013 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092605 pd=0.922174 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=5930,268
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2730,149
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.220489 ps=2.195652 w=1 l=0.15
**devattr s=5930,268 d=11000,510
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.092605 ps=0.922174 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.118032 ps=1.313948 w=0.65 l=0.15
**devattr s=4010,197 d=7150,370
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.564 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6600,266
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.07602 pd=0.866 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4872,284
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.07602 pd=0.866 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.182 ps=1.564 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07602 ps=0.866 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07602 pd=0.866 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=2814,151
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.564 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=12000,520
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07602 ps=0.866 w=0.42 l=0.15
**devattr s=2814,151 d=2352,140
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.182 ps=1.564 w=1 l=0.15
**devattr s=6600,266 d=5600,256
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.564 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR VNB VPB A X B_N
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.114071 ps=0.949948 w=0.42 l=0.15
**devattr s=6300,234 d=2268,138
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.114071 pd=0.949948 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=6300,234
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092605 pd=0.922174 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5930,268
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.176538 ps=1.470157 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.220489 ps=2.195652 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.092605 ps=0.922174 w=0.42 l=0.15
**devattr s=4368,272 d=4704,280
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114071 pd=0.949948 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.252686 pd=2.194215 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=12600,526
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.127562 pd=1.32793 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7410,374
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.252686 ps=2.194215 w=1 l=0.15
**devattr s=5930,268 d=5400,254
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.127562 ps=1.32793 w=0.65 l=0.15
**devattr s=4075,198 d=3510,184
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.082425 pd=0.858047 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.082425 ps=0.858047 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.082425 pd=0.858047 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.106128 pd=0.92157 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
.ends

.subckt sky130_fd_sc_hd__nor4_1 VPB VNB VGND VPWR Y D C B A
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.103188 pd=0.9675 as=0.129187 ps=1.3725 w=0.65 l=0.15
**devattr s=3575,185 d=3510,184
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
**devattr s=5200,252 d=7600,276
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.129187 pd=1.3725 as=0.103188 ps=0.9675 w=0.65 l=0.15
**devattr s=4745,203 d=3575,185
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.129187 pd=1.3725 as=0.103188 ps=0.9675 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
**devattr s=7600,276 d=5400,254
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5200,252
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.103188 pd=0.9675 as=0.129187 ps=1.3725 w=0.65 l=0.15
**devattr s=6760,364 d=4745,203
.ends

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196667 pd=1.726667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=6600,266
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.196667 ps=1.726667 w=1 l=0.15
**devattr s=6600,266 d=10400,504
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=6760,364
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.196667 ps=1.726667 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=10600,506
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
**devattr s=6200,262 d=10600,506
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.180375 pd=1.205 as=0.118083 ps=1.23 w=0.65 l=0.15
**devattr s=3640,186 d=4030,192
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.180375 pd=1.205 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=10400,290
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.180375 ps=1.205 w=0.65 l=0.15
**devattr s=10400,290 d=3640,186
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=3640,186
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=6200,262
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.180375 ps=1.205 w=0.65 l=0.15
**devattr s=4030,192 d=6890,366
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.076853 ps=0.850815 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.076853 ps=0.850815 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.087697 pd=0.792676 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.118939 ps=1.316738 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.208803 ps=1.887324 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.076853 pd=0.850815 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.076853 pd=0.850815 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
.ends

.subckt sky130_fd_sc_hd__nand4_2 VNB VPB VGND VPWR D C Y B A
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25625 pd=1.7625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=8600,286
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.147875 pd=1.43 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25625 ps=1.7625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25625 pd=1.7625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25625 pd=1.7625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=16800,568
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.131625 pd=1.38 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.131625 pd=1.38 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7280,372
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25625 ps=1.7625 w=1 l=0.15
**devattr s=13400,334 d=5400,254
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.147875 ps=1.43 w=0.65 l=0.15
**devattr s=7280,372 d=3510,184
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25625 pd=1.7625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=13400,334
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.147875 ps=1.43 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.131625 ps=1.38 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25625 ps=1.7625 w=1 l=0.15
**devattr s=8600,286 d=5400,254
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.147875 pd=1.43 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=9360,404
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25625 ps=1.7625 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.131625 ps=1.38 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.191667 ps=1.716667 w=1 l=0.15
**devattr s=6300,263 d=10400,504
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.104813 ps=0.9725 w=0.65 l=0.15
**devattr s=4095,193 d=6760,364
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.104813 ps=0.9725 w=0.65 l=0.15
**devattr s=4290,196 d=2730,172
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.191667 pd=1.716667 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6600,266 d=6300,263
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.191667 ps=1.716667 w=1 l=0.15
**devattr s=10400,504 d=6600,266
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=6760,364
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104813 pd=0.9725 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104813 pd=0.9725 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4095,193
.ends

.subckt sky130_fd_sc_hd__nor3_1 VPB VNB VGND VPWR C B A Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VNB VPB VPWR VGND X A1_N A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.128382 ps=1.053134 w=0.42 l=0.15
**devattr s=5830,267 d=5160,236
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=4368,272
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06831 pd=0.73445 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
**devattr s=2688,148 d=1764,126
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.06831 ps=0.73445 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128382 pd=1.053134 as=0.129 ps=1.18 w=0.42 l=0.15
**devattr s=5160,236 d=8370,269
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.128382 ps=1.053134 w=0.42 l=0.15
**devattr s=8370,269 d=2688,148
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.06831 ps=0.73445 w=0.42 l=0.15
**devattr s=3945,196 d=2646,147
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305672 pd=2.507463 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5830,267
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128382 pd=1.053134 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4368,272
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.105719 pd=1.136649 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3945,196
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VPB VNB VGND VPWR A1 A2 Y B2 C1 B1
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.113633 pd=1.22 as=0.14205 ps=1.415 w=0.65 l=0.15
**devattr s=6608,364 d=3510,184
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243333 pd=1.82 as=0.12 ps=1.24 w=1 l=0.15
**devattr s=4800,248 d=9000,290
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.013333 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14205 pd=1.415 as=0.113633 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=4680,202
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.34 ps=2.013333 w=1 l=0.15
**devattr s=15200,352 d=4800,248
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.243333 ps=1.82 w=1 l=0.15
**devattr s=9000,290 d=4200,242
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.013333 as=0.243333 ps=1.82 w=1 l=0.15
**devattr s=11200,512 d=15200,352
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.14205 ps=1.415 w=0.65 l=0.15
**devattr s=4680,202 d=3510,184
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14205 pd=1.415 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.113633 pd=1.22 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6616,364
.ends

.subckt sky130_fd_sc_hd__o221a_1 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=7280,372
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.388333 pd=2.11 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=16500,365
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.122417 pd=1.243333 as=0.2015 ps=1.92 w=0.65 l=0.15
**devattr s=8060,384 d=3965,191
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.122417 ps=1.243333 w=0.65 l=0.15
**devattr s=3965,191 d=3510,184
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6600,266
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=11200,512
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.122417 pd=1.243333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.388333 ps=2.11 w=1 l=0.15
**devattr s=13600,536 d=6600,266
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.388333 ps=2.11 w=1 l=0.15
**devattr s=16500,365 d=4200,242
.ends

.subckt sky130_fd_sc_hd__a221oi_1 VGND VPWR VPB VNB Y B1 C1 A1 A2 B2
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3965,191
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.14375 ps=1.2875 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14375 pd=1.2875 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.069875 pd=0.865 as=0.1365 ps=1.286667 w=0.65 l=0.15
**devattr s=4225,195 d=2795,173
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.286667 as=0.099125 ps=0.955 w=0.65 l=0.15
**devattr s=3965,191 d=7930,382
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14375 pd=1.2875 as=0.2825 ps=2.565 w=1 l=0.15
**devattr s=10400,504 d=6100,261
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.069875 ps=0.865 w=0.65 l=0.15
**devattr s=2795,173 d=6760,364
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2825 pd=2.565 as=0.14375 ps=1.2875 w=1 l=0.15
**devattr s=6100,261 d=12200,522
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.286667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4225,195
.ends

.subckt sky130_fd_sc_hd__o41a_1 VPB VNB VGND VPWR X B1 A4 A3 A2 A1
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1339 pd=1.192 as=0.1248 ps=1.164 w=0.65 l=0.15
**devattr s=3510,184 d=4940,206
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1248 pd=1.164 as=0.1339 ps=1.192 w=0.65 l=0.15
**devattr s=4940,206 d=5070,208
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.183333 ps=1.7 w=1 l=0.15
**devattr s=5400,254 d=10400,304
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.183333 pd=1.7 as=0.425 ps=2.85 w=1 l=0.15
**devattr s=17000,570 d=5400,254
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.1339 pd=1.192 as=0.247 ps=2.06 w=0.65 l=0.15
**devattr s=9880,412 d=6760,364
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1339 pd=1.192 as=0.1248 ps=1.164 w=0.65 l=0.15
**devattr s=5070,208 d=5070,208
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1248 pd=1.164 as=0.1339 ps=1.192 w=0.65 l=0.15
**devattr s=5070,208 d=7800,380
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
**devattr s=8800,288 d=7800,278
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=7800,278
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1248 pd=1.164 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
**devattr s=10400,304 d=8800,288
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.183333 pd=1.7 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=11200,512
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20625 pd=1.9125 as=0.16875 ps=1.5875 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091542 pd=0.931667 as=0.117 ps=1.226667 w=0.65 l=0.15
**devattr s=7280,372 d=3510,184
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.226667 as=0.091542 ps=0.931667 w=0.65 l=0.15
**devattr s=3965,191 d=6760,364
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14375 pd=1.2875 as=0.2025 ps=1.905 w=1 l=0.15
**devattr s=5400,254 d=6100,261
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.226667 as=0.134062 ps=1.3875 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.091542 ps=0.931667 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2025 pd=1.905 as=0.14375 ps=1.2875 w=1 l=0.15
**devattr s=6100,261 d=10400,504
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.226667 as=0.091542 ps=0.931667 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.134062 pd=1.3875 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.134062 ps=1.3875 w=0.65 l=0.15
**devattr s=7150,370 d=3510,184
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.134062 pd=1.3875 as=0.117 ps=1.226667 w=0.65 l=0.15
**devattr s=3510,184 d=7280,372
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.5875 as=0.20625 ps=1.9125 w=1 l=0.15
**devattr s=11000,510 d=5400,254
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2025 pd=1.905 as=0.16875 ps=1.5875 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.091542 pd=0.931667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.5875 as=0.2025 ps=1.905 w=1 l=0.15
**devattr s=11200,512 d=5400,254
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14375 pd=1.2875 as=0.16875 ps=1.5875 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.5875 as=0.14375 ps=1.2875 w=1 l=0.15
**devattr s=5400,254 d=11200,512
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091542 pd=0.931667 as=0.117 ps=1.226667 w=0.65 l=0.15
**devattr s=3510,184 d=3965,191
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20625 pd=1.9125 as=0.16875 ps=1.5875 w=1 l=0.15
**devattr s=5400,254 d=11200,512
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.5875 as=0.20625 ps=1.9125 w=1 l=0.15
**devattr s=5400,254 d=5400,254
.ends

.subckt sky130_fd_sc_hd__or4bb_1 VPWR VGND VPB VNB B A X D_N C_N
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.072904 pd=0.814826 as=0.058275 ps=0.6975 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.100675 pd=0.988673 as=0.05985 ps=0.705 w=0.42 l=0.15
**devattr s=2394,141 d=5930,268
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4860,266
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.072904 pd=0.814826 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2478,143
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.100675 pd=0.988673 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4904,264
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.239701 ps=2.353982 w=1 l=0.15
**devattr s=5930,268 d=11000,510
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.072904 pd=0.814826 as=0.058275 ps=0.6975 w=0.42 l=0.15
**devattr s=2394,141 d=2268,138
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2394,141
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.072904 ps=0.814826 w=0.42 l=0.15
**devattr s=2478,143 d=4368,272
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.100675 ps=0.988673 w=0.42 l=0.15
**devattr s=4904,264 d=4704,280
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
**devattr s=4860,266 d=1764,126
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.058275 pd=0.6975 as=0.072904 ps=0.814826 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.058275 pd=0.6975 as=0.072904 ps=0.814826 w=0.42 l=0.15
**devattr s=4368,272 d=2394,141
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.112827 ps=1.261041 w=0.65 l=0.15
**devattr s=4075,198 d=7150,370
.ends

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
**devattr s=2990,176 d=6760,364
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=12000,520
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=2730,172
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.2015 ps=1.92 w=0.65 l=0.15
**devattr s=6760,364 d=2990,176
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=9360,404
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.2925 ps=2.443662 w=1 l=0.15
**devattr s=6662,278 d=7800,278
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2925 pd=2.443662 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=15200,552
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.026338 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.114914 pd=1.01093 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.177843 ps=1.564535 w=0.65 l=0.15
**devattr s=4472,208 d=5070,208
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.177843 pd=1.564535 as=0.12675 ps=1.04 w=0.65 l=0.15
**devattr s=5070,208 d=9880,412
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12285 ps=1.026338 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.52 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.52 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.104 ps=1.1 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.104 ps=1.1 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.1 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.1 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.52 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.1 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4452,274
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.913333 as=0.083052 ps=0.789823 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.083052 ps=0.789823 w=0.42 l=0.15
**devattr s=6670,287 d=1764,126
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.083052 pd=0.789823 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.913333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112949 ps=1.025665 w=0.42 l=0.15
**devattr s=5544,216 d=2268,138
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112949 pd=1.025665 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112949 pd=1.025665 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=5544,216
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112949 ps=1.025665 w=0.42 l=0.15
**devattr s=4804,217 d=2268,138
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.197743 pd=1.880531 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=6670,287
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.174803 pd=1.587339 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4804,217
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
**devattr s=5850,220 d=5720,218
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.193 ps=1.586 w=1 l=0.15
**devattr s=7400,274 d=5600,256
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
**devattr s=5720,218 d=2730,172
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23375 pd=1.4675 as=0.33 ps=2.66 w=1 l=0.15
**devattr s=13200,532 d=9700,297
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.386667 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=6890,366
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.386667 w=0.65 l=0.15
**devattr s=6695,233 d=3900,190
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.586 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.386667 as=0.2145 ps=1.96 w=0.65 l=0.15
**devattr s=8580,392 d=6695,233
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.586 as=0.23375 ps=1.4675 w=1 l=0.15
**devattr s=9700,297 d=6600,266
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23375 pd=1.4675 as=0.193 ps=1.586 w=1 l=0.15
**devattr s=6600,266 d=9000,290
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.586 as=0.23375 ps=1.4675 w=1 l=0.15
**devattr s=9000,290 d=7400,274
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
**devattr s=3900,190 d=5850,220
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207025 pd=2.021472 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.207025 ps=2.021472 w=1 l=0.15
**devattr s=6030,269 d=5400,254
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.849018 as=0.085983 ps=0.996667 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.166109 pd=1.534302 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7150,370
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2142,135
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.849018 as=0.085983 ps=0.996667 w=0.42 l=0.15
**devattr s=2975,163 d=6030,269
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.166109 ps=1.534302 w=0.65 l=0.15
**devattr s=5216,221 d=3510,184
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.085983 pd=0.996667 as=0.08695 ps=0.849018 w=0.42 l=0.15
**devattr s=2268,138 d=2975,163
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.107332 pd=0.991395 as=0.05355 ps=0.675 w=0.42 l=0.15
**devattr s=2142,135 d=5216,221
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPB VNB VPWR VGND A1 B1_N Y A2
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
**devattr s=6100,261 d=5100,251
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06952 ps=0.781395 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4030,192
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.10759 ps=1.209302 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.263017 pd=2.214876 as=0.1275 ps=1.255 w=1 l=0.15
**devattr s=5100,251 d=11200,512
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10759 pd=1.209302 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=4030,192 d=3510,184
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.110467 pd=0.930248 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=7130,280
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.263017 ps=2.214876 w=1 l=0.15
**devattr s=7130,280 d=6100,261
.ends

.subckt sky130_fd_sc_hd__and4bb_1 VNB VPB VGND VPWR A_N B_N C D X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08715 pd=0.868636 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=3108,158 d=6880,292
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.081493 ps=0.796021 w=0.42 l=0.15
**devattr s=2352,140 d=5544,300
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2940,154
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.08715 ps=0.868636 w=0.42 l=0.15
**devattr s=2352,140 d=5376,296
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08715 pd=0.868636 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=6720,328 d=2352,140
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.081493 pd=0.796021 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=6720,328 d=2352,140
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=2.068182 w=1 l=0.15
**devattr s=6880,292 d=10400,504
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2352,140
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.081493 pd=0.796021 as=0.0777 ps=0.79 w=0.42 l=0.15
**devattr s=3108,158 d=5060,222
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.08715 ps=0.868636 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.08715 ps=0.868636 w=0.42 l=0.15
**devattr s=4872,284 d=2352,140
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.12612 ps=1.231937 w=0.65 l=0.15
**devattr s=5060,222 d=6616,364
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08715 pd=0.868636 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2352,140 d=2940,154
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20125 pd=1.9025 as=0.144167 ps=1.288333 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.129594 ps=1.37375 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.221667 pd=2.11 as=0.144167 ps=1.288333 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.144167 pd=1.288333 as=0.221667 ps=2.11 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.129594 ps=1.37375 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.096688 ps=0.9475 w=0.65 l=0.15
**devattr s=4225,195 d=6760,364
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.129594 pd=1.37375 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.129594 ps=1.37375 w=0.65 l=0.15
**devattr s=7150,370 d=3510,184
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.129594 pd=1.37375 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.144167 pd=1.288333 as=0.20125 ps=1.9025 w=1 l=0.15
**devattr s=11000,510 d=5400,254
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.221667 pd=2.11 as=0.144167 ps=1.288333 w=1 l=0.15
**devattr s=6500,265 d=10400,504
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.096688 pd=0.9475 as=0.129594 ps=1.37375 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.144167 pd=1.288333 as=0.221667 ps=2.11 w=1 l=0.15
**devattr s=5400,254 d=6500,265
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.129594 pd=1.37375 as=0.096688 ps=0.9475 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.129594 pd=1.37375 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20125 pd=1.9025 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.221667 ps=2.11 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.221667 pd=2.11 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=11200,512
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.096688 pd=0.9475 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=4225,195
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20125 ps=1.9025 w=1 l=0.15
**devattr s=5400,254 d=5400,254
.ends

.subckt sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21125 pd=1.9225 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.21125 ps=1.9225 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.41 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=4420,198
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.21125 ps=1.9225 w=1 l=0.15
**devattr s=6300,263 d=10400,504
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.141375 ps=1.41 w=0.65 l=0.15
**devattr s=6890,366 d=3640,186
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.141375 ps=1.41 w=0.65 l=0.15
**devattr s=4420,198 d=6500,230
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
**devattr s=6500,230 d=4940,206
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21125 pd=1.9225 as=0.18 ps=1.693333 w=1 l=0.15
**devattr s=5600,256 d=6300,263
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.41 as=0.1235 ps=1.03 w=0.65 l=0.15
**devattr s=4940,206 d=6890,366
.ends

.subckt top clk rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] uo_out[0] uo_out[1] uo_out[2]
+ uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VPWR VGND
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0985_ game.h\[0\] clknet_3_2__leaf_clk _0036_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0770_ VPWR VGND VGND VPWR _0295_ _0131_ _0313_ _0322_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0968_ game.ballY\[5\] clknet_3_1__leaf_clk _0019_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0899_ VGND VPWR _0435_ game.paddle\[6\] game.paddle\[7\] game.paddle\[8\] VPWR VGND
+ sky130_fd_sc_hd__and3_1
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ VGND VPWR _0369_ _0355_ _0372_ _0371_ _0364_ VPWR VGND sky130_fd_sc_hd__and4b_1
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ VGND VPWR _0027_ _0307_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0684_ VPWR VGND _0248_ game.ballY\[4\] _0244_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_19_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_147 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0805_ VPWR VGND VPWR VGND _0353_ _0351_ _0352_ _0355_ _0354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0598_ VGND VPWR _0006_ _0173_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0667_ _0233_ _0225_ game.ballY\[2\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0736_ VPWR VGND _0292_ game.ballX\[4\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_46_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0521_ VGND VPWR _0104_ _0105_ _0066_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1004_ game.v\[8\] clknet_3_4__leaf_clk _0055_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ VPWR VGND _0278_ _0277_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_37_17 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0504_ VPWR VGND VPWR VGND new_game.d net3 sky130_fd_sc_hd__inv_2
XFILLER_0_40_270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ game.inBallY clknet_3_4__leaf_clk _0035_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0967_ game.ballY\[4\] clknet_3_5__leaf_clk _0018_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0898_ VGND VPWR VPWR VGND _0434_ _0338_ _0339_ _0337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xmax_cap6 VGND VPWR net6 _0152_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0752_ VPWR VGND VGND VPWR _0307_ _0209_ _0306_ sky130_fd_sc_hd__or2_1
X_0821_ _0371_ _0357_ _0347_ _0356_ _0370_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ VPWR VGND VGND VPWR _0244_ game.ballY\[4\] _0247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0804_ VPWR VGND VGND VPWR _0065_ _0354_ game.ballX\[1\] sky130_fd_sc_hd__nand2_1
X_0735_ VGND VPWR _0025_ _0291_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0597_ VPWR VGND _0173_ _0172_ _0161_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0666_ _0232_ game.ballY\[2\] _0225_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0520_ VPWR VGND VPWR VGND _0102_ _0095_ _0103_ _0104_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ game.v\[7\] clknet_3_4__leaf_clk _0054_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0718_ VPWR VGND VPWR VGND _0276_ game.ballX\[1\] _0222_ _0277_ _0147_ sky130_fd_sc_hd__a22o_1
X_0649_ VGND VPWR _0216_ _0217_ _0168_ _0218_ _0208_ game.paddle\[8\] VPWR VGND sky130_fd_sc_hd__a41o_1
XFILLER_0_35_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0503_ VPWR VGND VPWR VGND pause.d net2 sky130_fd_sc_hd__inv_2
XFILLER_0_27_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0983_ game.ballDirX clknet_3_1__leaf_clk _0034_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0897_ VGND VPWR _0340_ _0433_ _0432_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0966_ game.ballY\[3\] clknet_3_5__leaf_clk _0017_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0751_ VPWR VGND VGND VPWR _0305_ _0257_ game.ballX\[5\] _0304_ _0306_ sky130_fd_sc_hd__o22a_1
X_0820_ VGND VPWR _0292_ _0370_ _0063_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0682_ VPWR VGND _0246_ _0239_ _0234_ _0231_ _0245_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_34_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0949_ game.paddle\[6\] clknet_3_4__leaf_clk _0011_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_0803_ VPWR VGND VGND VPWR _0353_ _0065_ game.ballX\[1\] sky130_fd_sc_hd__or2_1
X_0665_ VGND VPWR _0230_ _0221_ _0231_ _0226_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_0734_ VPWR VGND _0291_ _0290_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0596_ VGND VPWR VPWR VGND _0172_ _0171_ game.paddle\[1\] _0168_ sky130_fd_sc_hd__mux2_1
Xhold10 net16 game.inPaddle VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ game.v\[6\] clknet_3_1__leaf_clk _0053_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0648_ VGND VPWR _0211_ _0174_ _0217_ game.paddle\[7\] VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0717_ VGND VPWR _0275_ _0276_ game.ballX\[0\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0579_ VGND VPWR _0158_ game.offset\[2\] game.offset\[3\] _0150_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_35_214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0502_ VPWR VGND VPWR VGND game.h\[7\] _0089_ _0090_ game.hsync game.h\[9\] sky130_fd_sc_hd__nand4_1
XFILLER_0_27_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ game.ballDirY clknet_3_1__leaf_clk _0033_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0896_ VPWR VGND VGND VPWR game.paddle\[7\] _0432_ game.paddle\[6\] sky130_fd_sc_hd__nand2_1
X_0965_ game.ballY\[2\] clknet_3_5__leaf_clk _0016_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0750_ VPWR VGND VPWR VGND _0303_ _0302_ _0212_ _0305_ sky130_fd_sc_hd__a21o_1
X_0681_ VPWR VGND VGND VPWR game.ballY\[2\] game.ballY\[3\] _0244_ _0245_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0948_ game.paddle\[5\] clknet_3_5__leaf_clk _0010_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_0879_ VGND VPWR _0140_ _0410_ _0421_ _0066_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ VPWR VGND VGND VPWR _0064_ _0352_ game.ballX\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0664_ VPWR VGND VGND VPWR _0225_ _0230_ game.ballY\[1\] sky130_fd_sc_hd__nand2_1
X_0733_ VPWR VGND VPWR VGND _0289_ game.ballX\[3\] _0222_ _0290_ _0145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0595_ VPWR VGND VGND VPWR _0163_ _0167_ game.new_game_n _0171_ sky130_fd_sc_hd__o21a_1
Xhold11 net17 game.paddle\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ game.v\[5\] clknet_3_3__leaf_clk _0052_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0578_ VGND VPWR _0002_ _0157_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0647_ VPWR VGND _0216_ _0195_ game.paddle\[6\] game.paddle\[7\] _0174_ VGND VPWR
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0716_ VGND VPWR game.ballX\[1\] _0275_ game.ballDirX VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0501_ VPWR VGND VPWR VGND _0079_ _0066_ game.h\[8\] _0090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0981_ game.inBallX clknet_3_1__leaf_clk _0032_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0964_ game.ballY\[1\] clknet_3_5__leaf_clk _0015_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_0895_ VPWR VGND VPWR VGND _0428_ net11 _0431_ _0045_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0680_ VPWR VGND VPWR VGND _0244_ _0225_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0947_ game.paddle\[4\] clknet_3_7__leaf_clk _0009_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_0878_ VPWR VGND _0420_ _0140_ _0066_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0801_ VPWR VGND VGND VPWR _0351_ _0064_ game.ballX\[0\] sky130_fd_sc_hd__or2_1
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0594_ VGND VPWR _0005_ _0170_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0663_ VGND VPWR _0015_ _0229_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0732_ VGND VPWR _0288_ _0289_ _0287_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold12 net18 game.v\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1000_ game.v\[4\] clknet_3_6__leaf_clk _0051_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0715_ VGND VPWR VGND VPWR _0022_ _0273_ _0223_ _0274_ _0161_ sky130_fd_sc_hd__o211a_1
X_0577_ VGND VPWR _0157_ _0155_ _0138_ _0156_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0646_ VPWR VGND VGND VPWR _0209_ _0215_ _0012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0500_ VPWR VGND VPWR VGND _0066_ game.h\[6\] _0063_ _0089_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0629_ VGND VPWR _0197_ _0200_ _0201_ _0196_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0980_ game.hit clknet_3_3__leaf_clk _0031_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0894_ VGND VPWR _0428_ _0410_ _0431_ net11 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0963_ game.ballY\[0\] clknet_3_5__leaf_clk _0014_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_98 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0877_ VGND VPWR _0039_ _0419_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0946_ game.paddle\[3\] clknet_3_7__leaf_clk _0008_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0731_ VPWR VGND VPWR VGND _0283_ _0280_ _0282_ _0288_ sky130_fd_sc_hd__a21oi_1
X_0800_ VPWR VGND VPWR VGND _0346_ game.ballX\[7\] _0349_ _0350_ sky130_fd_sc_hd__a21oi_1
X_0593_ VGND VPWR _0170_ _0138_ net19 _0169_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0662_ VPWR VGND _0229_ _0228_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0929_ VGND VPWR _0457_ game.v\[6\] game.v\[7\] _0453_ VPWR VGND sky130_fd_sc_hd__and3_1
Xhold13 net19 game.paddle\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0645_ VGND VPWR VPWR VGND _0215_ _0210_ _0214_ game.paddle\[7\] sky130_fd_sc_hd__mux2_1
X_0714_ VPWR VGND VGND VPWR _0273_ _0274_ _0212_ sky130_fd_sc_hd__nand2_1
X_0576_ VPWR VGND VGND VPWR game.offset\[2\] _0156_ _0150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ VGND VPWR VGND VPWR _0200_ _0199_ _0198_ _0175_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0559_ game.h\[7\] game.h\[9\] _0141_ game.h\[8\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0962_ up_key.dff1 clknet_3_6__leaf_clk up_key.d VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0893_ VGND VPWR _0044_ _0430_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0945_ game.paddle\[2\] clknet_3_7__leaf_clk _0007_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0876_ _0140_ _0418_ _0419_ net1 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ VGND VPWR game.ballX\[3\] _0287_ game.ballDirX VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0661_ VPWR VGND VPWR VGND _0227_ game.ballY\[1\] _0223_ _0228_ _0147_ sky130_fd_sc_hd__a22o_1
X_0592_ VPWR VGND VGND VPWR _0169_ game.new_game_n _0168_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ VPWR VGND VPWR VGND _0396_ _0397_ _0392_ _0406_ _0405_ sky130_fd_sc_hd__or4b_1
XFILLER_0_30_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0928_ VGND VPWR VGND VPWR _0456_ net20 _0453_ _0053_ sky130_fd_sc_hd__o21ba_1
Xhold14 net20 game.v\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_215 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0644_ VPWR VGND VPWR VGND _0167_ _0214_ _0213_ _0174_ _0211_ _0212_ sky130_fd_sc_hd__a2111o_1
X_0713_ VPWR VGND VPWR VGND _0273_ game.ballX\[0\] sky130_fd_sc_hd__inv_2
X_0575_ VPWR VGND VGND VPWR _0155_ game.offset\[2\] _0150_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0558_ VGND VPWR VGND VPWR _0140_ game.h\[2\] game.h\[3\] game.h\[0\] game.h\[1\]
+ sky130_fd_sc_hd__and4_2
X_0627_ VGND VPWR _0181_ game.paddle\[5\] _0199_ game.paddle\[4\] VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0489_ VPWR VGND VPWR VGND game.v\[8\] _0057_ game.v\[9\] _0081_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ game.up_key_n clknet_3_7__leaf_clk net7 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0892_ _0428_ _0410_ _0430_ _0429_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_5_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0944_ game.paddle\[1\] clknet_3_7__leaf_clk _0006_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ VPWR VGND _0418_ _0065_ _0062_ _0064_ game.h\[3\] VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0591_ VPWR VGND VGND VPWR _0167_ _0168_ _0163_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0660_ VGND VPWR _0226_ _0227_ game.ballY\[0\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ VPWR VGND _0456_ _0450_ _0084_ game.v\[6\] _0209_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0789_ VGND VPWR VPWR VGND game.v\[8\] _0340_ game.paddle\[8\] sky130_fd_sc_hd__xor2_1
X_0858_ VGND VPWR VGND VPWR _0405_ _0133_ _0394_ _0401_ _0404_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 net21 game.v\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0574_ VGND VPWR _0001_ _0154_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0643_ VPWR VGND VPWR VGND _0195_ game.paddle\[6\] _0174_ _0213_ sky130_fd_sc_hd__a21oi_1
X_0712_ VPWR VGND VPWR VGND _0272_ _0266_ _0209_ _0021_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk VGND VPWR VGND VPWR clk clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0626_ VPWR VGND VPWR VGND game.paddle\[5\] _0181_ game.paddle\[4\] _0198_ sky130_fd_sc_hd__or3_1
X_0557_ VPWR VGND VGND VPWR game.h\[5\] game.h\[6\] _0139_ sky130_fd_sc_hd__nor2_1
X_0488_ VGND VPWR _0079_ game.h\[9\] _0080_ _0068_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0609_ VGND VPWR VPWR VGND _0174_ _0183_ game.paddle\[3\] game.paddle\[2\] game.paddle\[1\]
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0960_ down_key.dff1 clknet_3_7__leaf_clk down_key.d VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0891_ VPWR VGND VGND VPWR _0429_ game.h\[8\] _0426_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_111 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0943_ game.paddle\[0\] clknet_3_7__leaf_clk _0005_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0874_ VGND VPWR _0038_ _0417_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0590_ VPWR VGND VGND VPWR _0164_ _0166_ _0167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ VGND VPWR _0404_ _0402_ game.inBallY _0403_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0926_ VGND VPWR _0052_ _0455_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0788_ VGND VPWR VPWR VGND game.v\[7\] _0339_ game.paddle\[7\] sky130_fd_sc_hd__xor2_1
XFILLER_0_23_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold16 net22 game.h\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ VGND VPWR VPWR VGND _0212_ _0271_ _0270_ _0272_ sky130_fd_sc_hd__or3b_1
X_0573_ _0150_ _0138_ _0154_ _0153_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_20_183 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0642_ VGND VPWR _0163_ _0212_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_0909_ _0441_ _0138_ _0443_ _0442_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_43_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0625_ VPWR VGND VGND VPWR game.paddle\[5\] _0194_ _0197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0556_ VPWR VGND _0138_ net1 VPWR VGND sky130_fd_sc_hd__buf_2
X_0487_ VPWR VGND _0079_ game.h\[6\] _0063_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0608_ VPWR VGND VGND VPWR _0180_ _0182_ _0181_ sky130_fd_sc_hd__nand2_1
X_0539_ _0123_ _0113_ _0106_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0890_ VGND VPWR _0428_ game.h\[8\] game.h\[7\] _0423_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0942_ game.offset\[4\] clknet_3_2__leaf_clk _0004_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0873_ VGND VPWR _0417_ _0415_ _0138_ _0416_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_50_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ VGND VPWR VGND VPWR game.v\[6\] _0338_ game.paddle\[6\] sky130_fd_sc_hd__or2b_1
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0856_ VGND VPWR VPWR VGND game.v\[4\] _0403_ game.ballY\[3\] sky130_fd_sc_hd__xor2_1
X_0925_ _0453_ net1 _0455_ _0454_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold17 net23 game.inBallX VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0641_ VPWR VGND VGND VPWR _0211_ game.paddle\[6\] _0198_ sky130_fd_sc_hd__or2_1
X_0710_ VPWR VGND VPWR VGND _0268_ _0267_ _0264_ _0271_ _0269_ sky130_fd_sc_hd__a22o_1
X_0572_ VPWR VGND _0153_ _0152_ game.pause_n game.offset\[0\] game.offset\[1\] VGND
+ VPWR sky130_fd_sc_hd__a31o_1
X_0908_ VPWR VGND VGND VPWR _0442_ game.v\[1\] _0438_ sky130_fd_sc_hd__or2_1
X_0839_ VGND VPWR VPWR VGND game.v\[7\] _0386_ game.ballY\[6\] sky130_fd_sc_hd__xor2_1
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0624_ VPWR VGND VGND VPWR _0196_ _0174_ _0195_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0555_ VPWR VGND VPWR VGND _0137_ _0084_ game.hit game.speaker game.v\[6\] sky130_fd_sc_hd__a22o_1
X_0486_ VGND VPWR _0078_ game.v\[7\] game.v\[8\] game.v\[6\] VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_202 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0538_ VGND VPWR _0121_ _0122_ _0102_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0607_ VGND VPWR VPWR VGND game.paddle\[2\] game.paddle\[1\] game.paddle\[3\] _0181_
+ sky130_fd_sc_hd__or3_2
X_0469_ VPWR VGND _0062_ game.h\[0\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_39_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ game.offset\[3\] clknet_3_2__leaf_clk _0003_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0872_ VPWR VGND VPWR VGND _0062_ _0064_ _0065_ _0416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0924_ VPWR VGND VGND VPWR _0454_ _0084_ _0450_ sky130_fd_sc_hd__or2_1
X_0786_ VGND VPWR VGND VPWR game.paddle\[6\] _0337_ game.v\[6\] sky130_fd_sc_hd__or2b_1
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0855_ VGND VPWR game.ballY\[2\] _0402_ game.v\[3\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0571_ VPWR VGND VGND VPWR _0152_ _0143_ _0151_ _0073_ _0058_ sky130_fd_sc_hd__nor4_1
X_0640_ VGND VPWR _0168_ game.paddle\[7\] _0210_ game.new_game_n VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0907_ VGND VPWR _0441_ game.v\[0\] game.v\[1\] _0142_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0769_ VPWR VGND VPWR VGND _0312_ _0317_ _0311_ _0321_ sky130_fd_sc_hd__or3_1
X_0838_ VPWR VGND VGND VPWR game.ballY\[6\] game.ballY\[7\] _0385_ _0384_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0623_ VPWR VGND _0195_ _0194_ game.paddle\[5\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0554_ VGND VPWR VGND VPWR _0137_ _0132_ _0134_ game.ballX\[8\] _0136_ sky130_fd_sc_hd__a211o_1
X_0485_ VPWR VGND VPWR VGND _0064_ _0065_ _0066_ _0077_ game.h\[3\] sky130_fd_sc_hd__nand4_1
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0537_ _0121_ _0103_ _0095_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0606_ VGND VPWR game.paddle\[1\] game.paddle\[3\] _0180_ game.paddle\[2\] VPWR VGND
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0468_ VPWR VGND VGND VPWR _0058_ _0061_ game.row0 sky130_fd_sc_hd__nor2_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_3_2__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ game.offset\[2\] clknet_3_2__leaf_clk _0002_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0871_ VPWR VGND VGND VPWR _0064_ _0062_ _0415_ _0065_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ VPWR VGND VPWR VGND _0399_ _0398_ _0400_ _0401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0923_ VPWR VGND _0453_ _0450_ _0084_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0785_ VPWR VGND VPWR VGND _0330_ _0335_ _0333_ _0151_ _0336_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0570_ VGND VPWR VGND VPWR _0141_ _0140_ _0151_ _0139_ game.h\[4\] sky130_fd_sc_hd__nand4_2
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0906_ VPWR VGND VGND VPWR _0438_ _0440_ _0047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0837_ VGND VPWR _0384_ game.ballY\[4\] game.ballY\[3\] game.ballY\[5\] VPWR VGND
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0768_ VPWR VGND VGND VPWR _0209_ _0320_ _0029_ sky130_fd_sc_hd__nor2_1
X_0699_ VGND VPWR game.ballY\[6\] _0261_ _0225_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0622_ _0194_ game.paddle\[2\] game.paddle\[4\] game.paddle\[3\] game.paddle\[1\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0484_ VPWR VGND VPWR VGND game.v\[4\] _0071_ _0076_ _0072_ _0073_ _0075_ sky130_fd_sc_hd__a221o_1
X_0553_ VPWR VGND VGND VPWR _0135_ game.ballY\[7\] game.ballY\[6\] _0136_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0536_ VGND VPWR _0119_ _0120_ _0109_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0605_ VGND VPWR _0007_ _0179_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0467_ VPWR VGND VPWR VGND game.v\[8\] _0060_ game.v\[3\] _0059_ _0061_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0519_ _0103_ game.offset\[4\] game.h\[3\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_36_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ VGND VPWR _0037_ _0414_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0999_ game.v\[3\] clknet_3_6__leaf_clk _0050_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0922_ VGND VPWR _0051_ _0452_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0853_ VGND VPWR VPWR VGND game.v\[1\] _0400_ game.ballY\[0\] sky130_fd_sc_hd__xor2_1
X_0784_ VPWR VGND VPWR VGND game.v\[3\] _0331_ _0335_ game.paddle\[1\] _0071_ _0334_
+ sky130_fd_sc_hd__a221o_1
Xinput1 VGND VPWR rst_n net1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0905_ VGND VPWR _0142_ _0439_ _0440_ net21 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0767_ VGND VPWR VPWR VGND _0320_ game.ballX\[7\] _0223_ _0319_ _0318_ sky130_fd_sc_hd__o2bb2a_1
X_0836_ VGND VPWR _0034_ _0383_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0698_ VGND VPWR _0260_ game.ballY\[6\] game.new_game_n _0212_ VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0621_ VPWR VGND _0193_ net1 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0483_ VPWR VGND VGND VPWR game.v\[4\] _0074_ _0075_ sky130_fd_sc_hd__nor2_1
X_0552_ VPWR VGND VGND VPWR _0135_ game.ballY\[4\] game.ballY\[5\] sky130_fd_sc_hd__or2_1
XFILLER_0_17_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ VPWR VGND VPWR VGND _0369_ _0359_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0604_ VGND VPWR _0179_ _0169_ _0138_ _0178_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0535_ VGND VPWR _0118_ _0119_ _0099_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0466_ VPWR VGND VPWR VGND game.v\[1\] game.v\[0\] game.v\[2\] _0060_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0518_ VGND VPWR _0100_ _0101_ _0102_ _0099_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0998_ game.v\[2\] clknet_3_6__leaf_clk _0049_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0921_ _0450_ _0138_ _0452_ _0451_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0783_ VGND VPWR VPWR VGND game.v\[4\] _0334_ game.paddle\[4\] sky130_fd_sc_hd__xor2_1
X_0852_ VPWR VGND VGND VPWR game.v\[2\] _0399_ game.ballY\[1\] sky130_fd_sc_hd__nand2_1
Xinput2 VGND VPWR net2 ui_in[0] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0904_ VPWR VGND VGND VPWR _0208_ net6 _0439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ VPWR VGND VPWR VGND _0343_ _0382_ _0209_ _0383_ sky130_fd_sc_hd__or3_1
X_0697_ VGND VPWR _0019_ _0259_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0766_ VPWR VGND _0319_ _0317_ _0315_ _0310_ _0212_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0620_ VGND VPWR _0009_ _0192_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0551_ VGND VPWR VGND VPWR _0134_ game.ballY\[5\] _0133_ game.ballY\[7\] game.ballY\[6\]
+ sky130_fd_sc_hd__o211a_1
X_0482_ VPWR VGND VPWR VGND _0074_ game.v\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_17_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_84 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0749_ VPWR VGND VGND VPWR _0302_ _0303_ _0304_ sky130_fd_sc_hd__nor2_1
X_0818_ VPWR VGND VPWR VGND _0350_ _0363_ _0348_ _0368_ _0367_ sky130_fd_sc_hd__or4b_1
X_0603_ VGND VPWR VPWR VGND _0178_ _0145_ _0177_ game.paddle\[2\] _0168_ sky130_fd_sc_hd__o2bb2a_1
X_0534_ VGND VPWR VPWR VGND game.v\[2\] _0118_ _0065_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0465_ VPWR VGND _0059_ game.v\[9\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0517_ VGND VPWR VGND VPWR game.offset\[3\] _0101_ _0065_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0997_ game.v\[1\] clknet_3_6__leaf_clk _0048_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0920_ VPWR VGND VGND VPWR _0451_ game.v\[4\] _0447_ sky130_fd_sc_hd__or2_1
X_0782_ VPWR VGND VGND VPWR game.v\[3\] _0331_ _0333_ _0071_ _0332_ game.paddle\[1\]
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_23_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0851_ VPWR VGND VGND VPWR _0398_ game.v\[2\] game.ballY\[1\] sky130_fd_sc_hd__or2_1
Xinput3 VGND VPWR net3 ui_in[1] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0903_ VPWR VGND _0438_ _0142_ game.v\[0\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_28_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0834_ VPWR VGND VGND VPWR _0381_ _0080_ _0295_ _0382_ sky130_fd_sc_hd__o21a_1
X_0765_ VPWR VGND VPWR VGND _0315_ _0310_ _0317_ _0318_ sky130_fd_sc_hd__a21oi_1
X_0696_ VPWR VGND VGND VPWR _0259_ _0209_ _0258_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_229 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0550_ VPWR VGND _0133_ game.ballY\[4\] game.ballY\[3\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0481_ VPWR VGND VGND VPWR game.v\[3\] _0073_ game.v\[2\] sky130_fd_sc_hd__nand2_1
X_0817_ VPWR VGND VGND VPWR _0365_ _0063_ _0359_ _0358_ _0367_ _0366_ sky130_fd_sc_hd__o221a_1
X_0679_ VGND VPWR _0017_ _0243_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0748_ VPWR VGND VPWR VGND _0298_ _0294_ _0297_ _0303_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0533_ VGND VPWR VPWR VGND _0117_ _0093_ _0116_ _0091_ _0092_ _0094_ sky130_fd_sc_hd__a221oi_1
X_0602_ VGND VPWR VPWR VGND _0177_ _0175_ _0176_ _0164_ sky130_fd_sc_hd__mux2_1
X_0464_ VPWR VGND VGND VPWR _0058_ game.v\[4\] _0057_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0516_ _0100_ _0065_ game.offset\[3\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_162 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_118 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0996_ game.v\[0\] clknet_3_6__leaf_clk _0047_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ VPWR VGND VGND VPWR _0059_ _0385_ _0397_ sky130_fd_sc_hd__nor2_1
X_0781_ VPWR VGND VGND VPWR _0087_ game.paddle\[5\] _0328_ game.paddle\[2\] _0332_
+ sky130_fd_sc_hd__o22a_1
Xinput4 VGND VPWR net4 ui_in[2] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ game.ballX\[8\] clknet_3_1__leaf_clk _0030_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0902_ VPWR VGND VGND VPWR _0342_ _0437_ _0161_ _0046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0833_ VPWR VGND VPWR VGND _0381_ game.inBallX sky130_fd_sc_hd__inv_2
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0695_ VGND VPWR VPWR VGND _0258_ _0255_ _0256_ game.ballY\[5\] _0257_ sky130_fd_sc_hd__o2bb2a_1
X_0764_ VGND VPWR VPWR VGND _0295_ _0317_ game.ballX\[7\] sky130_fd_sc_hd__xor2_1
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0480_ VPWR VGND VGND VPWR _0072_ game.v\[2\] game.v\[1\] sky130_fd_sc_hd__or2_1
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0747_ VGND VPWR VPWR VGND _0295_ _0302_ game.ballX\[5\] sky130_fd_sc_hd__xor2_1
X_0816_ VPWR VGND VPWR VGND _0292_ game.ballX\[3\] _0364_ _0366_ sky130_fd_sc_hd__a21o_1
X_0678_ VPWR VGND _0243_ _0242_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0601_ VGND VPWR VPWR VGND game.paddle\[2\] _0176_ game.paddle\[1\] sky130_fd_sc_hd__xor2_1
X_0532_ VGND VPWR _0115_ _0116_ _0105_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0463_ VPWR VGND VPWR VGND game.v\[6\] game.v\[5\] game.v\[7\] _0057_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0515_ VPWR VGND VPWR VGND _0097_ _0096_ _0098_ _0099_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0995_ game.inPaddle clknet_3_6__leaf_clk _0046_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0780_ VPWR VGND VPWR VGND _0331_ game.paddle\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_23_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput5 VGND VPWR net5 ui_in[3] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ game.ballX\[7\] clknet_3_0__leaf_clk _0029_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_206 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0901_ VPWR VGND VGND VPWR _0437_ net16 _0436_ _0434_ _0433_ _0336_ sky130_fd_sc_hd__o41a_1
X_0763_ VPWR VGND VPWR VGND _0316_ _0308_ _0209_ _0028_ sky130_fd_sc_hd__a21oi_1
X_0832_ VPWR VGND VPWR VGND _0380_ _0378_ _0209_ _0033_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0694_ VPWR VGND VGND VPWR game.new_game_n _0257_ _0212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0746_ VGND VPWR _0026_ _0301_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0815_ VPWR VGND VGND VPWR _0130_ _0365_ _0364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0677_ VPWR VGND VPWR VGND _0241_ game.ballY\[3\] _0223_ _0242_ _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0531_ VGND VPWR _0114_ _0115_ game.v\[4\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0600_ VPWR VGND _0175_ _0166_ _0174_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0729_ VGND VPWR _0024_ _0286_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0514_ _0098_ game.offset\[2\] _0064_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_35_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0994_ game.h\[9\] clknet_3_2__leaf_clk _0045_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0977_ game.ballX\[6\] clknet_3_1__leaf_clk _0028_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0900_ VGND VPWR VPWR VGND _0059_ _0436_ _0435_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0762_ VGND VPWR VPWR VGND _0314_ _0315_ _0212_ _0316_ sky130_fd_sc_hd__or3b_1
X_0693_ VPWR VGND VGND VPWR _0256_ _0253_ _0254_ sky130_fd_sc_hd__or2_1
X_0831_ VGND VPWR _0081_ _0244_ _0380_ _0379_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0814_ VGND VPWR game.ballX\[5\] _0364_ game.h\[6\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0676_ VGND VPWR _0240_ _0241_ _0239_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0745_ VPWR VGND _0301_ _0300_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0530_ VPWR VGND VPWR VGND _0112_ _0106_ _0113_ _0114_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1013_ VGND VPWR game.row0 uo_out[7] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ VPWR VGND _0286_ _0285_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0659_ VGND VPWR _0226_ _0225_ game.ballY\[1\] VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0513_ VGND VPWR VGND VPWR _0062_ _0097_ game.offset\[1\] sky130_fd_sc_hd__or2b_1
XFILLER_0_39_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0993_ game.h\[8\] clknet_3_2__leaf_clk _0044_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0976_ game.ballX\[5\] clknet_3_0__leaf_clk _0027_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0830_ VPWR VGND VPWR VGND _0379_ game.inBallY sky130_fd_sc_hd__inv_2
XFILLER_0_11_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0692_ VPWR VGND VPWR VGND _0254_ _0253_ _0212_ _0255_ sky130_fd_sc_hd__a21oi_1
X_0761_ VPWR VGND VPWR VGND _0313_ _0312_ _0311_ _0315_ sky130_fd_sc_hd__a21o_1
X_0959_ down_key.dff2 clknet_3_7__leaf_clk net8 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ VPWR VGND VPWR VGND _0356_ _0355_ _0363_ _0362_ _0357_ sky130_fd_sc_hd__or4bb_1
X_0675_ VPWR VGND VPWR VGND _0234_ _0231_ _0233_ _0240_ sky130_fd_sc_hd__a21oi_1
X_0744_ VPWR VGND VPWR VGND _0299_ _0292_ _0222_ _0300_ _0145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ VGND VPWR game.col0 uo_out[6] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0727_ VPWR VGND VPWR VGND _0284_ game.ballX\[2\] _0222_ _0285_ _0145_ sky130_fd_sc_hd__a22o_1
X_0589_ VPWR VGND VGND VPWR _0166_ _0165_ game.paddle\[8\] game.paddle\[5\] game.paddle\[6\]
+ game.paddle\[7\] sky130_fd_sc_hd__o41a_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0658_ VGND VPWR game.ballDirY _0225_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0512_ VGND VPWR VGND VPWR game.h\[1\] _0096_ game.offset\[2\] sky130_fd_sc_hd__or2b_1
XFILLER_0_39_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0992_ game.h\[7\] clknet_3_0__leaf_clk _0043_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0975_ game.ballX\[4\] clknet_3_0__leaf_clk _0026_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0760_ VGND VPWR _0314_ _0312_ _0311_ _0313_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0691_ VGND VPWR game.ballY\[5\] _0254_ _0225_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0958_ new_game.dff1 clknet_3_7__leaf_clk new_game.d VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0889_ VPWR VGND VGND VPWR _0426_ _0427_ _0043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ VGND VPWR VPWR VGND _0294_ _0299_ _0298_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0812_ VPWR VGND VPWR VGND _0063_ _0361_ _0362_ _0358_ _0359_ sky130_fd_sc_hd__a22oi_1
X_0674_ VPWR VGND VPWR VGND _0239_ _0238_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1011_ VGND VPWR game.speaker uo_out[5] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0726_ VGND VPWR VPWR VGND _0280_ _0284_ _0283_ sky130_fd_sc_hd__xor2_1
X_0588_ VPWR VGND VPWR VGND _0165_ game.up_key_n sky130_fd_sc_hd__inv_2
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0657_ VGND VPWR VGND VPWR _0014_ _0221_ _0223_ _0224_ _0161_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0511_ VGND VPWR VGND VPWR game.h\[3\] _0095_ game.offset\[4\] sky130_fd_sc_hd__or2b_1
XFILLER_0_39_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ _0270_ _0268_ _0267_ _0264_ _0269_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0991_ game.h\[6\] clknet_3_2__leaf_clk _0042_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ game.ballX\[3\] clknet_3_0__leaf_clk _0025_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0690_ VPWR VGND VPWR VGND _0249_ _0246_ _0248_ _0253_ sky130_fd_sc_hd__a21oi_1
X_0957_ game.new_game_n clknet_3_7__leaf_clk net9 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0888_ VGND VPWR _0423_ _0410_ _0427_ net22 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0673_ VGND VPWR VPWR VGND _0225_ _0238_ game.ballY\[3\] sky130_fd_sc_hd__xor2_1
X_0742_ VPWR VGND VGND VPWR _0296_ _0297_ _0298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0811_ VPWR VGND VGND VPWR _0130_ _0361_ _0360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1010_ VGND VPWR game.vsync uo_out[4] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_0725_ VPWR VGND VGND VPWR _0281_ _0282_ _0283_ sky130_fd_sc_hd__nor2_1
X_0656_ VPWR VGND VGND VPWR _0221_ _0224_ _0212_ sky130_fd_sc_hd__nand2_1
X_0587_ VPWR VGND VPWR VGND game.paddle\[8\] game.paddle\[7\] down_key.dff2 _0164_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0510_ VGND VPWR VGND VPWR game.v\[0\] _0094_ game.offset\[1\] sky130_fd_sc_hd__or2b_1
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 net7 up_key.dff1 VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0639_ VGND VPWR VGND VPWR _0011_ _0206_ _0207_ _0204_ _0209_ sky130_fd_sc_hd__a211o_1
X_0708_ VPWR VGND VGND VPWR _0225_ _0269_ game.ballY\[7\] sky130_fd_sc_hd__nand2_1
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ game.h\[5\] clknet_3_3__leaf_clk _0041_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0973_ game.ballX\[2\] clknet_3_0__leaf_clk _0024_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ pause.dff1 clknet_3_7__leaf_clk pause.d VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ VPWR VGND _0426_ _0423_ game.h\[7\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_33_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0810_ VPWR VGND VGND VPWR game.ballX\[3\] _0360_ _0292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0741_ _0297_ _0295_ _0292_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0672_ VGND VPWR _0016_ _0237_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0939_ game.offset\[1\] clknet_3_3__leaf_clk _0001_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0586_ VPWR VGND VGND VPWR _0163_ game.pause_n net6 sky130_fd_sc_hd__nand2_2
X_0655_ VGND VPWR _0222_ _0223_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_0724_ _0282_ game.ballDirX game.ballX\[2\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold2 net8 down_key.dff1 VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ VPWR VGND VGND VPWR _0268_ _0225_ game.ballY\[7\] sky130_fd_sc_hd__or2_1
XFILLER_0_29_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0569_ VGND VPWR _0150_ game.offset\[0\] game.offset\[1\] _0145_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0638_ VGND VPWR _0208_ _0209_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ game.ballX\[1\] clknet_3_0__leaf_clk _0023_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_161 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0955_ game.pause_n clknet_3_7__leaf_clk net10 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0886_ VGND VPWR _0042_ _0425_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0740_ _0296_ _0292_ _0295_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0671_ VPWR VGND _0237_ _0236_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0938_ game.offset\[0\] clknet_3_3__leaf_clk _0000_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0869_ VGND VPWR _0414_ _0410_ _0412_ _0413_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_30_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ _0281_ game.ballX\[2\] game.ballDirX VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0585_ VPWR VGND VPWR VGND _0158_ net12 _0162_ _0004_ sky130_fd_sc_hd__a21oi_1
X_0654_ VPWR VGND game.new_game_n _0222_ _0163_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_34_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 net9 new_game.dff1 VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0706_ VPWR VGND VGND VPWR _0244_ _0267_ game.ballY\[6\] sky130_fd_sc_hd__nand2_1
X_0568_ VGND VPWR _0000_ _0149_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0499_ VPWR VGND VGND VPWR _0078_ _0075_ game.vsync _0088_ sky130_fd_sc_hd__nand3_1
X_0637_ VPWR VGND VPWR VGND _0208_ net1 sky130_fd_sc_hd__inv_2
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0971_ game.ballX\[0\] clknet_3_0__leaf_clk _0022_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0954_ qb clknet_3_6__leaf_clk game.blue VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_224 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0885_ _0423_ _0410_ _0425_ _0424_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0670_ VPWR VGND VPWR VGND _0235_ game.ballY\[2\] _0223_ _0236_ _0147_ sky130_fd_sc_hd__a22o_1
X_0868_ VPWR VGND VGND VPWR _0413_ _0064_ _0062_ sky130_fd_sc_hd__or2_1
X_0937_ VPWR VGND VPWR VGND _0460_ _0059_ _0462_ _0056_ sky130_fd_sc_hd__a21oi_1
X_0799_ VGND VPWR game.ballX\[8\] _0349_ game.h\[9\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0722_ VGND VPWR _0279_ _0273_ _0280_ _0275_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_0653_ VPWR VGND VPWR VGND _0221_ game.ballY\[0\] sky130_fd_sc_hd__inv_2
X_0584_ VGND VPWR _0158_ _0161_ _0162_ net12 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold4 net10 pause.dff1 VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0636_ VPWR VGND VPWR VGND _0169_ _0204_ _0206_ _0207_ sky130_fd_sc_hd__a21oi_1
X_0705_ VPWR VGND VGND VPWR net13 _0266_ _0223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0498_ VGND VPWR _0087_ _0059_ _0088_ game.v\[1\] _0084_ VPWR VGND sky130_fd_sc_hd__and4b_1
X_0567_ VGND VPWR _0149_ _0146_ _0138_ _0148_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0619_ VPWR VGND _0192_ _0191_ _0161_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0970_ game.ballY\[7\] clknet_3_5__leaf_clk _0021_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ qg clknet_3_3__leaf_clk game.green VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0884_ VPWR VGND _0424_ _0140_ _0066_ _0063_ game.h\[6\] VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0936_ VGND VPWR _0460_ _0439_ _0462_ _0059_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ VPWR VGND VGND VPWR _0064_ _0412_ _0062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ VGND VPWR _0347_ _0348_ _0346_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0652_ VGND VPWR _0013_ _0220_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0583_ VPWR VGND _0161_ net1 VPWR VGND sky130_fd_sc_hd__buf_4
X_0721_ VPWR VGND VGND VPWR game.ballDirX _0279_ game.ballX\[1\] sky130_fd_sc_hd__nand2_1
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0919_ VGND VPWR _0450_ game.v\[3\] game.v\[4\] _0444_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 net11 game.h\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0566_ VPWR VGND VGND VPWR game.offset\[0\] _0148_ _0147_ sky130_fd_sc_hd__nand2_1
X_0635_ VGND VPWR _0206_ _0196_ _0168_ _0205_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_20_63 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0704_ VPWR VGND VGND VPWR _0260_ _0265_ _0161_ _0020_ sky130_fd_sc_hd__o21a_1
X_0497_ VPWR VGND VPWR VGND _0087_ game.v\[2\] sky130_fd_sc_hd__inv_2
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0618_ VPWR VGND VPWR VGND _0190_ game.paddle\[4\] _0171_ _0191_ _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0549_ VGND VPWR VGND VPWR _0132_ _0130_ game.ballX\[5\] _0131_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0952_ qr clknet_3_3__leaf_clk game.red VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ VGND VPWR _0423_ _0079_ _0066_ _0140_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_10_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0866_ VGND VPWR _0036_ _0411_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ VGND VPWR VGND VPWR _0055_ net18 _0457_ _0461_ _0161_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ VGND VPWR game.ballX\[7\] _0347_ game.h\[8\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ VGND VPWR _0023_ _0278_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0582_ VGND VPWR _0003_ _0160_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0651_ _0220_ _0218_ _0219_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0918_ VGND VPWR _0050_ _0449_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0849_ VPWR VGND VPWR VGND game.ballY\[3\] _0393_ _0396_ _0394_ _0133_ _0395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold6 net12 game.offset\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0703_ VGND VPWR _0265_ _0263_ _0147_ _0264_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0496_ VPWR VGND VPWR VGND _0086_ _0082_ _0085_ game.green sky130_fd_sc_hd__a21oi_1
X_0634_ VPWR VGND VGND VPWR _0174_ _0205_ _0198_ sky130_fd_sc_hd__nand2_1
X_0565_ VGND VPWR _0145_ _0147_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_195 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0479_ VPWR VGND VPWR VGND _0071_ game.v\[1\] sky130_fd_sc_hd__inv_2
X_0617_ VGND VPWR VGND VPWR _0189_ _0167_ _0188_ _0190_ game.paddle\[4\] sky130_fd_sc_hd__a2bb2o_1
X_0548_ VPWR VGND VGND VPWR game.ballX\[6\] game.ballX\[7\] _0131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0951_ game.paddle\[8\] clknet_3_5__leaf_clk _0013_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_0882_ VPWR VGND VPWR VGND _0420_ _0063_ _0422_ _0041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0865_ _0411_ _0062_ _0410_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0934_ VPWR VGND VPWR VGND _0461_ _0460_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0796_ _0346_ game.ballX\[5\] game.ballX\[3\] _0292_ game.ballX\[6\] VGND VPWR VPWR
+ VGND sky130_fd_sc_hd__and4_1
X_0581_ _0158_ _0138_ _0160_ _0159_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0650_ VGND VPWR VPWR VGND _0219_ _0217_ _0216_ _0168_ _0169_ game.paddle\[8\] sky130_fd_sc_hd__a32o_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0917_ _0447_ _0439_ _0449_ _0448_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0779_ VPWR VGND VPWR VGND _0328_ game.paddle\[5\] _0330_ game.paddle\[2\] _0087_
+ _0329_ sky130_fd_sc_hd__a221o_1
X_0848_ VGND VPWR _0393_ _0142_ _0395_ game.ballY\[3\] VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold7 net13 game.ballY\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0633_ VPWR VGND VPWR VGND _0204_ net17 sky130_fd_sc_hd__inv_2
X_0702_ VPWR VGND VGND VPWR _0261_ _0264_ _0262_ sky130_fd_sc_hd__nand2_1
X_0564_ VPWR VGND VGND VPWR _0146_ game.offset\[0\] _0145_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0495_ VPWR VGND VGND VPWR game.inBallY _0086_ net23 sky130_fd_sc_hd__nand2_1
XFILLER_0_9_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0616_ VPWR VGND _0189_ _0181_ _0166_ _0174_ _0183_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0478_ VGND VPWR VPWR VGND _0069_ game.inPaddle _0063_ _0070_ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0547_ VPWR VGND VGND VPWR _0130_ game.ballX\[3\] game.ballX\[4\] sky130_fd_sc_hd__or2_1
XFILLER_0_48_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0881_ VGND VPWR _0420_ _0410_ _0422_ _0063_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0950_ game.paddle\[7\] clknet_3_4__leaf_clk _0012_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_0795_ VGND VPWR _0031_ _0345_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0864_ VPWR VGND VGND VPWR _0142_ _0410_ _0208_ sky130_fd_sc_hd__nor2_2
X_0933_ VGND VPWR _0460_ _0078_ _0084_ _0450_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_2_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0580_ VPWR VGND VPWR VGND _0150_ game.offset\[2\] game.offset\[3\] _0159_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ VPWR VGND VGND VPWR _0448_ game.v\[3\] _0444_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ VGND VPWR VPWR VGND game.v\[0\] _0329_ game.paddle\[0\] sky130_fd_sc_hd__xor2_1
X_0847_ VGND VPWR game.ballY\[5\] _0394_ game.v\[6\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 net14 game.ballX\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0563_ _0142_ _0145_ game.pause_n _0144_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_0632_ VGND VPWR _0010_ _0203_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0701_ VPWR VGND VGND VPWR _0263_ _0261_ _0262_ sky130_fd_sc_hd__or2_1
X_0494_ VPWR VGND VPWR VGND _0083_ _0070_ _0085_ game.red sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0546_ VGND VPWR VGND VPWR game.blue _0117_ _0127_ _0128_ _0129_ sky130_fd_sc_hd__o211a_1
X_0615_ VGND VPWR VGND VPWR _0188_ _0181_ _0183_ _0174_ game.paddle\[4\] sky130_fd_sc_hd__a211o_1
XFILLER_0_40_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0477_ VPWR VGND VGND VPWR game.col0 _0069_ _0067_ _0063_ _0062_ sky130_fd_sc_hd__nor4_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0529_ VPWR VGND VGND VPWR _0074_ game.offset\[4\] _0113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ VPWR VGND VGND VPWR _0420_ _0421_ _0040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ VGND VPWR _0054_ _0459_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0794_ _0342_ _0344_ _0345_ net1 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0863_ VGND VPWR VGND VPWR _0035_ _0391_ _0406_ _0161_ _0409_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0915_ VGND VPWR _0447_ game.v\[2\] game.v\[3\] _0441_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0777_ VPWR VGND VPWR VGND _0328_ _0084_ sky130_fd_sc_hd__inv_2
X_0846_ VGND VPWR game.ballY\[4\] _0393_ _0084_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold9 net15 game.inBallY VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_151 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0700_ VGND VPWR VPWR VGND _0262_ _0254_ _0249_ _0246_ _0135_ _0244_ sky130_fd_sc_hd__a32o_1
X_0562_ VPWR VGND VGND VPWR _0143_ _0073_ _0058_ _0144_ sky130_fd_sc_hd__nor3_1
X_0631_ VPWR VGND _0203_ _0202_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0493_ VPWR VGND VPWR VGND game.h\[9\] _0068_ _0085_ _0078_ _0084_ _0059_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0829_ VGND VPWR _0078_ net15 _0378_ _0059_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0614_ VGND VPWR _0008_ _0187_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0545_ VGND VPWR VGND VPWR _0129_ _0085_ _0070_ _0082_ _0086_ sky130_fd_sc_hd__o211a_1
X_0476_ VPWR VGND VPWR VGND game.h\[9\] _0068_ game.h\[6\] _0069_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0528_ VPWR VGND VPWR VGND _0110_ _0109_ _0111_ _0112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0862_ VPWR VGND _0409_ _0408_ _0407_ _0142_ game.inBallY VGND VPWR sky130_fd_sc_hd__a31o_1
X_0931_ _0457_ net1 _0459_ _0458_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_48_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0793_ VPWR VGND VPWR VGND game.hit game.new_game_n _0343_ _0344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0914_ VGND VPWR _0049_ _0446_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ VPWR VGND VPWR VGND _0384_ game.ballY\[6\] _0389_ _0392_ sky130_fd_sc_hd__a21oi_1
X_0776_ VGND VPWR _0030_ _0327_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0561_ VPWR VGND VPWR VGND game.v\[1\] game.v\[0\] game.v\[8\] _0143_ game.v\[9\]
+ sky130_fd_sc_hd__or4b_1
X_0630_ VPWR VGND VPWR VGND _0201_ game.paddle\[5\] _0171_ _0202_ _0147_ sky130_fd_sc_hd__a22o_1
X_0492_ VGND VPWR game.v\[5\] _0084_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_0759_ VPWR VGND VPWR VGND _0292_ _0295_ _0313_ game.ballX\[5\] sky130_fd_sc_hd__o21bai_1
X_0828_ VGND VPWR _0032_ _0377_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0613_ VPWR VGND _0187_ _0186_ _0161_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0544_ VGND VPWR VGND VPWR _0116_ _0128_ _0126_ sky130_fd_sc_hd__or2b_1
X_0475_ VPWR VGND VGND VPWR _0068_ game.h\[7\] game.h\[8\] sky130_fd_sc_hd__or2_1
XFILLER_0_0_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0527_ VPWR VGND VGND VPWR _0087_ game.offset\[3\] _0111_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0792_ VPWR VGND VGND VPWR _0070_ _0086_ _0343_ sky130_fd_sc_hd__nor2_1
X_0861_ _0403_ _0401_ _0408_ _0389_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0930_ VPWR VGND _0458_ _0450_ _0084_ game.v\[6\] game.v\[7\] VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_23_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0913_ _0444_ _0439_ _0446_ _0445_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0775_ VPWR VGND _0327_ _0326_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0844_ VPWR VGND VPWR VGND _0059_ _0385_ _0391_ _0387_ _0388_ _0390_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0491_ VPWR VGND _0083_ _0077_ _0076_ _0067_ _0082_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0560_ VGND VPWR VGND VPWR _0142_ _0141_ _0140_ _0139_ game.h\[4\] sky130_fd_sc_hd__and4_2
XFILLER_0_43_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0758_ VPWR VGND VPWR VGND _0302_ _0297_ _0296_ _0312_ _0294_ sky130_fd_sc_hd__or4b_1
X_0827_ VGND VPWR _0377_ _0374_ _0138_ _0376_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0689_ VGND VPWR _0018_ _0252_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0612_ VPWR VGND VPWR VGND _0185_ game.paddle\[3\] _0171_ _0186_ _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0543_ _0127_ _0092_ _0116_ _0091_ _0126_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0474_ VPWR VGND VPWR VGND game.h\[3\] _0066_ _0065_ _0064_ _0067_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0526_ VPWR VGND VGND VPWR _0087_ _0110_ game.offset\[3\] sky130_fd_sc_hd__nand2_1
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ VPWR VGND uo_out[3] game.hsync VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0509_ VGND VPWR VGND VPWR game.offset\[1\] _0093_ game.v\[0\] sky130_fd_sc_hd__or2b_1
XFILLER_0_17_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ VGND VPWR _0338_ _0336_ _0342_ _0341_ _0337_ VPWR VGND sky130_fd_sc_hd__and4b_1
XFILLER_0_23_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ VGND VPWR _0394_ _0386_ _0407_ _0402_ _0393_ VPWR VGND sky130_fd_sc_hd__and4b_1
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ game.h\[4\] clknet_3_3__leaf_clk _0040_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ VPWR VGND VGND VPWR _0445_ game.v\[2\] _0441_ sky130_fd_sc_hd__or2_1
X_0774_ VGND VPWR VGND VPWR game.ballX\[8\] _0324_ _0325_ _0326_ _0223_ sky130_fd_sc_hd__a2bb2o_1
X_0843_ VGND VPWR _0390_ _0389_ game.ballY\[6\] _0384_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0490_ VGND VPWR VGND VPWR _0059_ _0078_ _0080_ _0081_ _0082_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_29_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0757_ VPWR VGND VGND VPWR _0309_ _0311_ _0310_ sky130_fd_sc_hd__nand2_1
X_0688_ VPWR VGND _0252_ _0251_ _0193_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0826_ VPWR VGND VGND VPWR game.ballX\[8\] _0376_ _0375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0542_ VGND VPWR _0125_ _0126_ _0120_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0611_ VPWR VGND VPWR VGND _0183_ _0175_ _0182_ _0185_ _0184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0473_ VPWR VGND _0066_ game.h\[4\] VPWR VGND sky130_fd_sc_hd__buf_2
X_0809_ VPWR VGND _0359_ game.ballX\[6\] game.h\[7\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_31_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0525_ VPWR VGND VPWR VGND _0094_ _0107_ _0108_ _0109_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1008_ VPWR VGND uo_out[2] qr VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_44_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0508_ VPWR VGND VGND VPWR game.v\[0\] _0092_ _0062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0790_ VPWR VGND VGND VPWR _0339_ _0340_ _0341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ game.h\[3\] clknet_3_2__leaf_clk _0039_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0911_ VPWR VGND _0444_ _0441_ game.v\[2\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0842_ VGND VPWR game.ballY\[7\] _0389_ game.v\[8\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ VPWR VGND _0325_ _0323_ _0322_ _0321_ _0163_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_24_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ VGND VPWR VGND VPWR _0375_ game.ballX\[5\] game.ballX\[6\] _0292_ game.ballX\[7\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0756_ VGND VPWR VGND VPWR _0295_ _0310_ game.ballX\[6\] sky130_fd_sc_hd__or2b_1
X_0687_ VPWR VGND VPWR VGND _0250_ game.ballY\[4\] _0223_ _0251_ _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0541_ VGND VPWR VPWR VGND _0122_ _0125_ _0124_ sky130_fd_sc_hd__xor2_1
X_0610_ VPWR VGND VPWR VGND game.paddle\[1\] game.paddle\[2\] game.paddle\[3\] _0184_
+ sky130_fd_sc_hd__a21o_1
X_0472_ VPWR VGND _0065_ game.h\[2\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0808_ VPWR VGND VGND VPWR game.ballX\[3\] _0292_ _0358_ game.ballX\[5\] sky130_fd_sc_hd__nand3_1
X_0739_ VGND VPWR game.ballDirX _0295_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0524_ _0108_ game.offset\[2\] game.v\[1\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_1007_ VGND VPWR qg uo_out[1] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XPHY_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0507_ VPWR VGND VGND VPWR _0091_ game.v\[0\] _0062_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ game.h\[2\] clknet_3_2__leaf_clk _0038_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ VGND VPWR _0048_ _0443_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0772_ VPWR VGND VPWR VGND _0322_ _0321_ _0323_ _0324_ sky130_fd_sc_hd__a21oi_1
X_0841_ VPWR VGND VGND VPWR _0386_ _0388_ _0384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0755_ VGND VPWR VGND VPWR game.ballX\[6\] _0309_ _0295_ sky130_fd_sc_hd__or2b_1
X_0824_ VPWR VGND VPWR VGND _0373_ game.inBallX _0368_ _0374_ _0349_ sky130_fd_sc_hd__a22o_1
X_0686_ VGND VPWR VPWR VGND _0246_ _0250_ _0249_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_3_0__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0540_ VGND VPWR _0123_ _0124_ _0112_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0471_ VPWR VGND _0064_ game.h\[1\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0738_ VPWR VGND _0294_ _0287_ _0283_ _0280_ _0293_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0807_ VGND VPWR game.ballX\[2\] _0357_ game.h\[3\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0669_ VGND VPWR VPWR VGND _0231_ _0235_ _0234_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0523_ VGND VPWR VGND VPWR game.v\[1\] _0107_ game.offset\[2\] sky130_fd_sc_hd__or2b_1
X_1006_ VGND VPWR qb uo_out[0] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XPHY_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_268 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0506_ VPWR VGND VPWR VGND up_key.d net5 sky130_fd_sc_hd__inv_2
XFILLER_0_41_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ game.h\[1\] clknet_3_2__leaf_clk _0037_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_16 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0771_ VGND VPWR VPWR VGND _0295_ _0323_ game.ballX\[8\] sky130_fd_sc_hd__xor2_1
X_0840_ VPWR VGND VGND VPWR _0387_ _0386_ _0384_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ game.ballY\[6\] clknet_3_1__leaf_clk _0020_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0754_ VPWR VGND VGND VPWR net14 _0308_ _0223_ sky130_fd_sc_hd__nand2_1
X_0685_ VPWR VGND VGND VPWR _0247_ _0248_ _0249_ sky130_fd_sc_hd__nor2_1
X_0823_ VPWR VGND _0373_ _0346_ game.ballX\[7\] game.inBallX _0372_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_27_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0470_ VPWR VGND _0063_ game.h\[5\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_0_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0668_ VPWR VGND VGND VPWR _0232_ _0233_ _0234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0737_ VGND VPWR VGND VPWR game.ballDirX game.ballX\[2\] game.ballX\[3\] _0293_ sky130_fd_sc_hd__o21ba_1
X_0806_ VGND VPWR game.ballX\[3\] _0356_ _0066_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0599_ VGND VPWR VGND VPWR game.paddle\[8\] game.paddle\[7\] down_key.dff2 _0174_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_39_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0522_ VPWR VGND VGND VPWR _0074_ _0106_ game.offset\[4\] sky130_fd_sc_hd__nand2_1
XFILLER_0_21_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ game.v\[9\] clknet_3_4__leaf_clk _0056_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0505_ VPWR VGND VPWR VGND down_key.d net4 sky130_fd_sc_hd__inv_2
.ends

.subckt tt_um_argunda_tiny_opamp clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VPWR VGND
Xvbias_resistor_0 VPWR opamp_1/VBIAS VGND vbias_resistor
Xopamp_0 opamp_1/VBIAS VPWR ua[2] ua[1] ua[0] VGND opamp
Xopamp_1 opamp_1/VBIAS VPWR ua[5] ua[4] ua[3] VGND opamp
Xtop_0 clk rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] uo_out[0] uo_out[1] uo_out[2]
+ uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VPWR VGND top
R0 VGND uio_out[5] 0.000000
R1 VGND uio_out[6] 0.000000
R2 VGND uio_out[7] 0.000000
R3 VGND uio_oe[0] 0.000000
R4 VGND uio_oe[1] 0.000000
R5 VGND uio_oe[3] 0.000000
R6 VGND uio_oe[2] 0.000000
R7 VGND uio_out[0] 0.000000
R8 VGND uio_oe[4] 0.000000
R9 VGND uio_out[1] 0.000000
R10 VGND uio_out[2] 0.000000
R11 VGND uio_oe[5] 0.000000
R12 VGND uio_oe[6] 0.000000
R13 VGND uio_out[3] 0.000000
R14 VGND uio_oe[7] 0.000000
R15 VGND uio_out[4] 0.000000
.ends

