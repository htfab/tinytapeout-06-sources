magic
tech sky130A
magscale 1 2
timestamp 1713553032
<< nwell >>
rect -200 2630 990 2640
rect 360 1400 430 2630
<< pwell >>
rect 1140 2040 1800 2100
rect 1140 1380 1240 2040
rect 1680 1380 1800 2040
rect 1140 1300 1800 1380
rect 1140 1280 2000 1300
rect -400 1120 2000 1280
rect -400 480 -300 1120
rect 120 480 260 1120
rect 420 540 620 1080
rect 700 480 840 1120
rect 1280 480 1420 1120
rect 1840 480 2000 1120
rect -400 200 2000 480
<< psubdiff >>
rect 1700 1300 1800 2100
rect 1380 1220 1800 1240
rect -340 1140 1880 1220
rect 1380 1130 1880 1140
rect 1380 1120 1420 1130
rect 1830 1120 1880 1130
rect 1400 1090 1420 1120
<< locali >>
rect -400 2700 2000 2800
rect -400 2450 -340 2700
rect -360 1520 -340 2450
rect -220 2580 -180 2700
rect 940 2580 1060 2700
rect -220 2568 -68 2580
rect 260 2568 532 2580
rect 860 2568 1060 2580
rect -220 2540 1060 2568
rect -220 2506 -120 2540
rect -220 1532 -164 2506
rect -130 1532 -120 2506
rect 300 2506 480 2540
rect 300 2380 322 2506
rect 242 1650 322 2380
rect -220 1520 -120 1532
rect -360 1480 -120 1520
rect 300 1532 322 1650
rect 356 1532 436 2506
rect 470 2380 480 2506
rect 900 2520 1060 2540
rect 1860 2520 2000 2700
rect 900 2506 2000 2520
rect 780 2466 830 2480
rect 720 2407 830 2466
rect 470 1650 550 2380
rect 470 1532 480 1650
rect 720 1631 808 2407
rect 720 1572 830 1631
rect 780 1550 830 1572
rect 300 1480 480 1532
rect 900 1532 922 2506
rect 956 2450 2000 2506
rect 956 2176 1786 2450
rect 956 1532 1020 2176
rect 900 1480 1020 1532
rect -360 1470 1020 1480
rect -360 1436 -68 1470
rect 260 1436 532 1470
rect 860 1436 1020 1470
rect -360 1420 1020 1436
rect 1140 2040 1800 2100
rect 1140 2020 1240 2040
rect 1140 1320 1160 2020
rect 1220 1380 1240 2020
rect 1680 2020 1800 2040
rect 1680 1380 1700 2020
rect 1220 1360 1700 1380
rect 1220 1326 1292 1360
rect 1620 1326 1700 1360
rect 1220 1320 1700 1326
rect 1760 1320 1800 2020
rect 1140 1300 1800 1320
rect -400 1260 2000 1300
rect -400 1150 -340 1260
rect -400 1140 140 1150
rect 1860 1140 2000 1260
rect -400 1120 2000 1140
rect -400 1088 -300 1120
rect -400 532 -364 1088
rect -330 920 -300 1088
rect 120 1090 260 1120
rect -160 998 40 1080
rect -330 620 -220 920
rect -160 622 8 998
rect -330 532 -300 620
rect -160 560 40 622
rect -40 540 40 560
rect -400 480 -300 532
rect 120 530 150 1090
rect 250 920 260 1090
rect 700 1090 840 1120
rect 420 998 620 1080
rect 250 620 360 920
rect 420 622 588 998
rect 250 530 260 620
rect 420 540 620 622
rect 120 480 260 530
rect 700 530 720 1090
rect 820 920 840 1090
rect 1300 1090 1420 1120
rect 820 620 960 920
rect 820 530 840 620
rect 1170 610 1230 1010
rect 700 480 840 530
rect 1300 530 1310 1090
rect 1410 920 1420 1090
rect 1840 1088 2000 1120
rect 1410 622 1490 920
rect 1524 622 1540 920
rect 1410 620 1540 622
rect 1410 530 1420 620
rect 1300 490 1420 530
rect 1290 480 1420 490
rect 1840 532 1862 1088
rect 1896 532 2000 1088
rect 1840 480 2000 532
rect -400 440 2000 480
rect -400 300 -300 440
rect 1900 300 2000 440
rect -400 200 2000 300
<< viali >>
rect -340 1520 -220 2700
rect -180 2580 940 2700
rect -68 2568 260 2580
rect 532 2568 860 2580
rect -164 1532 -130 2506
rect 208 1631 242 2407
rect 322 1532 356 2506
rect 436 1532 470 2506
rect 1060 2520 1860 2700
rect 612 2466 780 2500
rect 550 1631 584 2407
rect 808 1631 842 2407
rect 612 1538 780 1572
rect 922 1532 956 2506
rect -68 1436 260 1470
rect 532 1436 860 1470
rect 1160 1320 1220 2020
rect 1372 1938 1540 1972
rect 1372 1428 1540 1462
rect 1292 1326 1620 1360
rect 1700 1320 1760 2020
rect -340 1150 1860 1260
rect 140 1140 1860 1150
rect -364 532 -330 1088
rect 8 622 42 998
rect 150 530 250 1090
rect 588 622 622 998
rect 720 530 820 1090
rect 1310 530 1410 1090
rect 1552 1048 1720 1082
rect 1490 622 1524 998
rect 1552 538 1720 572
rect 1862 532 1896 1088
rect -300 300 1900 440
<< metal1 >>
rect -400 2700 2000 2800
rect -400 2450 -340 2700
rect -360 1520 -340 2450
rect -220 2580 -180 2700
rect 940 2580 1060 2700
rect -220 2568 -68 2580
rect 260 2568 532 2580
rect 860 2568 1060 2580
rect -220 2540 1060 2568
rect -220 2506 -120 2540
rect -220 1532 -164 2506
rect -130 1532 -120 2506
rect 220 2506 560 2540
rect 40 2440 160 2500
rect 60 2280 160 2440
rect 220 2407 322 2506
rect 30 2220 40 2280
rect 140 2220 160 2280
rect -90 1660 -80 2020
rect 0 1660 10 2020
rect 60 1580 160 2220
rect 242 1631 322 2407
rect 220 1620 322 1631
rect 40 1560 160 1580
rect 40 1540 140 1560
rect -220 1520 -120 1532
rect -360 1480 -120 1520
rect 240 1532 322 1620
rect 356 1532 436 2506
rect 470 2407 560 2506
rect 906 2520 1060 2540
rect 1860 2520 2000 2700
rect 906 2506 2000 2520
rect 780 2466 840 2500
rect 620 2407 840 2466
rect 470 1631 550 2407
rect 620 2280 808 2407
rect 620 2220 680 2280
rect 760 2220 808 2280
rect 620 1631 808 2220
rect 470 1532 560 1631
rect 620 1620 840 1631
rect 620 1578 680 1620
rect 600 1572 680 1578
rect 760 1572 840 1620
rect 600 1538 612 1572
rect 780 1540 840 1572
rect 780 1538 792 1540
rect 600 1532 792 1538
rect 906 1532 922 2506
rect 956 2450 2000 2506
rect 956 2176 1786 2450
rect 956 1532 1020 2176
rect 240 1480 560 1532
rect 906 1484 1020 1532
rect 900 1480 1020 1484
rect -360 1470 1020 1480
rect -360 1436 -68 1470
rect 260 1436 532 1470
rect 860 1436 1020 1470
rect -360 1420 1020 1436
rect 1140 2040 1800 2100
rect 1140 2020 1240 2040
rect 1140 1320 1160 2020
rect 1220 1380 1240 2020
rect 1680 2020 1800 2040
rect 1370 1978 1380 1980
rect 1360 1972 1380 1978
rect 1520 1978 1530 1980
rect 1520 1972 1552 1978
rect 1360 1938 1372 1972
rect 1540 1938 1552 1972
rect 1360 1932 1380 1938
rect 1370 1920 1380 1932
rect 1520 1932 1552 1938
rect 1520 1920 1530 1932
rect 1380 1900 1520 1920
rect 1270 1810 1360 1840
rect 1270 1530 1280 1810
rect 1340 1530 1360 1810
rect 1270 1520 1360 1530
rect 1270 1510 1350 1520
rect 1410 1500 1500 1900
rect 1530 1830 1640 1860
rect 1530 1590 1550 1830
rect 1620 1590 1640 1830
rect 1530 1550 1640 1590
rect 1550 1500 1640 1550
rect 1410 1490 1520 1500
rect 1380 1468 1520 1490
rect 1360 1462 1552 1468
rect 1360 1428 1372 1462
rect 1540 1428 1552 1462
rect 1360 1422 1552 1428
rect 1380 1420 1520 1422
rect 1680 1380 1700 2020
rect 1220 1360 1700 1380
rect 1220 1326 1292 1360
rect 1620 1326 1700 1360
rect 1220 1320 1700 1326
rect 1760 1320 1800 2020
rect 1140 1300 1800 1320
rect 1140 1280 2000 1300
rect -400 1260 2000 1280
rect -400 1150 -340 1260
rect -400 1140 140 1150
rect 1860 1140 2000 1260
rect -400 1088 -300 1140
rect 120 1120 2000 1140
rect -400 532 -364 1088
rect -330 920 -300 1088
rect -198 1048 -188 1100
rect 20 1080 30 1100
rect 120 1090 260 1120
rect -170 1020 -160 1048
rect 20 1020 40 1080
rect -160 998 40 1020
rect -330 620 -220 920
rect -160 820 8 998
rect -160 760 -120 820
rect -60 760 8 820
rect -160 622 8 760
rect -330 532 -300 620
rect -160 560 40 622
rect -40 540 40 560
rect -400 480 -300 532
rect 120 530 150 1090
rect 250 920 260 1090
rect 700 1090 840 1120
rect 420 998 620 1080
rect 250 620 360 920
rect 420 820 588 998
rect 420 760 460 820
rect 520 760 588 820
rect 420 622 588 760
rect 250 530 260 620
rect 420 540 620 622
rect 120 480 260 530
rect 700 530 720 1090
rect 820 920 840 1090
rect 1300 1090 1420 1120
rect 1840 1110 2000 1120
rect 820 620 960 920
rect 1000 820 1120 1080
rect 1000 760 1040 820
rect 1100 760 1120 820
rect 820 530 840 620
rect 1000 540 1120 760
rect 1170 1000 1260 1010
rect 1170 900 1180 1000
rect 1260 900 1270 1000
rect 1170 610 1260 900
rect 700 480 840 530
rect 1300 530 1310 1090
rect 1410 920 1420 1090
rect 1850 1088 2000 1110
rect 1410 622 1490 920
rect 1524 622 1540 920
rect 1410 620 1540 622
rect 1580 830 1700 1048
rect 1580 770 1610 830
rect 1670 770 1700 830
rect 1410 530 1420 620
rect 1580 572 1700 770
rect 1750 840 1810 1000
rect 1750 610 1810 730
rect 1300 490 1420 530
rect 1290 480 1420 490
rect 1850 532 1862 1088
rect 1896 532 2000 1088
rect 1850 480 2000 532
rect -400 440 2000 480
rect -400 300 -300 440
rect 1900 300 2000 440
rect -400 200 2000 300
<< via1 >>
rect 40 2220 140 2280
rect -80 1660 0 2020
rect 680 2220 760 2280
rect 680 1572 760 1620
rect 680 1540 760 1572
rect 1380 1972 1520 1980
rect 1380 1938 1520 1972
rect 1380 1920 1520 1938
rect 1280 1530 1340 1810
rect 1550 1590 1620 1830
rect -188 1048 20 1100
rect -160 1020 20 1048
rect -120 760 -60 820
rect 460 760 520 820
rect 1040 760 1100 820
rect 1180 900 1260 1000
rect 1610 770 1670 830
rect 1750 730 1810 840
<< metal2 >>
rect -400 2300 -200 2360
rect 1800 2300 2000 2360
rect -400 2280 160 2300
rect -400 2220 40 2280
rect 140 2220 160 2280
rect -400 2200 160 2220
rect 640 2280 2000 2300
rect 640 2220 680 2280
rect 760 2220 2000 2280
rect 640 2200 2000 2220
rect -400 2160 -200 2200
rect -160 2020 80 2100
rect -160 1660 -80 2020
rect 0 1660 80 2020
rect -160 1260 80 1660
rect -200 1100 80 1260
rect 660 1620 780 2200
rect 1800 2160 2000 2200
rect 1380 1980 1520 1990
rect 1380 1910 1520 1920
rect 660 1540 680 1620
rect 760 1540 780 1620
rect 660 1230 780 1540
rect 1240 1810 1360 1860
rect 1240 1530 1280 1810
rect 1340 1530 1360 1810
rect 1550 1830 1620 1840
rect 1620 1590 2000 1760
rect 1550 1580 2000 1590
rect 1240 1380 1360 1530
rect 1560 1500 2000 1580
rect 1240 1280 1820 1380
rect 660 1130 1280 1230
rect -200 1048 -188 1100
rect -200 1020 -160 1048
rect 20 1020 80 1100
rect -200 980 80 1020
rect 1160 1000 1280 1130
rect -140 840 -20 980
rect 440 840 560 980
rect 1000 840 1120 1000
rect 1160 900 1180 1000
rect 1260 900 1280 1000
rect 1160 870 1280 900
rect 1730 840 1820 1280
rect -140 830 1700 840
rect -140 820 1610 830
rect -140 760 -120 820
rect -60 760 460 820
rect 520 760 1040 820
rect 1100 770 1610 820
rect 1670 770 1700 830
rect 1100 760 1700 770
rect -140 600 -20 760
rect 440 580 560 760
rect 1000 580 1120 760
rect 1730 730 1750 840
rect 1810 730 1820 840
rect 1730 720 1820 730
<< metal3 >>
rect 1380 2700 1520 2800
rect 1400 2100 1500 2700
rect 1300 1900 1600 2100
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM1
timestamp 1713470961
transform 1 0 96 0 1 2019
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM2
timestamp 1713470961
transform 1 0 696 0 1 2019
box -296 -619 296 619
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM3
timestamp 1713539272
transform 1 0 -104 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM4
timestamp 1713539272
transform 1 0 476 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM5
timestamp 1713539272
transform 1 0 1056 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM6
timestamp 1713539272
transform 1 0 1636 0 1 810
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM7
timestamp 1713539272
transform 1 0 1456 0 1 1700
box -296 -410 296 410
<< labels >>
flabel metal1 -400 2700 -300 2800 0 FreeSans 1600 0 0 0 VDD
port 4 nsew
flabel metal2 1836 2188 1970 2326 0 FreeSans 1600 0 0 0 VREF_OUT
port 6 nsew
flabel metal2 -378 2186 -244 2324 0 FreeSans 1600 0 0 0 VREF_IN
port 0 nsew
flabel pwell -392 204 -162 438 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel metal3 1380 2700 1520 2800 0 FreeSans 1600 0 0 0 OE
port 2 nsew
flabel metal2 1820 1550 1960 1710 0 FreeSans 1600 0 0 0 IOUT
port 3 nsew
<< end >>
