magic
tech sky130A
magscale 1 2
timestamp 1713422843
<< psubdiff >>
rect 1988 -2658 2060 -2118
rect 2078 -2658 3382 -2650
rect 1988 -2674 3382 -2658
rect 2060 -2684 3382 -2674
rect 2078 -2700 3382 -2684
<< locali >>
rect 1988 2830 7988 2900
rect 1988 2642 2240 2830
rect 1988 1628 2028 2642
rect 7920 2526 7988 2830
rect 3122 2398 4426 2526
rect 3122 1628 3242 2398
rect 1988 -566 3242 1628
rect 4312 2052 4426 2398
rect 6488 2406 7988 2526
rect 6488 2052 6606 2406
rect 6860 2404 7988 2406
rect 4312 1152 6606 2052
rect 4312 -566 5382 1152
rect 1988 -624 5382 -566
rect 1988 -626 5352 -624
rect 1988 -1568 3394 -730
rect 4160 -1568 5570 -730
rect 6286 -942 6596 1152
rect 7128 -914 7988 2404
rect 7124 -942 7988 -914
rect 6286 -1048 7988 -942
rect 1988 -2124 5578 -1568
rect 1988 -2658 2060 -2124
rect 2066 -2130 5578 -2124
rect 4112 -2136 5570 -2130
rect 4096 -2472 5574 -2136
rect 6092 -2456 7988 -1240
rect 6100 -2472 7988 -2456
rect 4096 -2516 7988 -2472
rect 4096 -2566 5128 -2516
rect 4118 -2616 5128 -2566
rect 4086 -2632 5128 -2616
rect 3980 -2648 5128 -2632
rect 3300 -2650 5128 -2648
rect 2078 -2658 5128 -2650
rect 1988 -2736 5128 -2658
rect 7906 -2736 7988 -2516
rect 1988 -3040 2228 -2736
rect 7908 -3040 7988 -2736
rect 1988 -3096 7988 -3040
rect 1988 -3100 7878 -3096
<< viali >>
rect 2240 2642 7920 2830
rect 2028 2526 7920 2642
rect 2028 1628 3122 2526
rect 4426 2052 6488 2526
rect 5128 -2736 7906 -2516
rect 2228 -3040 7908 -2736
<< metal1 >>
rect 1988 2830 7988 2900
rect 1988 2642 2240 2830
rect 1988 1628 2028 2642
rect 7920 2526 7988 2830
rect 3122 2482 4426 2526
rect 3122 1628 3178 2482
rect 3326 2344 3702 2482
rect 3326 2322 3420 2344
rect 3402 2272 3420 2322
rect 3608 2322 3702 2344
rect 3860 2354 4236 2482
rect 3608 2272 3626 2322
rect 3860 2312 3956 2354
rect 3946 2274 3956 2312
rect 4138 2312 4236 2354
rect 4138 2274 4148 2312
rect 3328 2220 3374 2244
rect 3662 2242 3898 2268
rect 3328 2218 3376 2220
rect 1988 -110 3178 1628
rect 3326 2088 3376 2218
rect 3658 2088 3898 2242
rect 3326 2052 4232 2088
rect 4362 2052 4426 2482
rect 6488 2484 7222 2526
rect 6488 2052 6576 2484
rect 6682 2389 7056 2435
rect 7210 2392 7222 2484
rect 6682 2213 6728 2389
rect 6762 2246 6772 2342
rect 6970 2246 6980 2342
rect 7010 2214 7056 2389
rect 3326 2036 3376 2052
rect 3326 1888 3370 2036
rect 3658 1894 3898 2052
rect 4362 1952 6576 2052
rect 6686 1906 6724 2213
rect 6762 2090 6772 2186
rect 6970 2090 6980 2186
rect 6760 1930 6770 2026
rect 6968 1930 6978 2026
rect 6632 1896 6724 1906
rect 3326 1860 3374 1888
rect 3656 1860 3898 1894
rect 6598 1876 6724 1896
rect 3326 1814 3898 1860
rect 3326 1792 3374 1814
rect 3656 1800 3898 1814
rect 3326 1654 3370 1792
rect 3658 1654 3898 1800
rect 3936 1796 3946 1870
rect 4148 1796 4158 1870
rect 6518 1788 6528 1876
rect 6666 1788 6724 1876
rect 6598 1756 6724 1788
rect 6760 1774 6770 1870
rect 6968 1774 6978 1870
rect 3326 1618 4222 1654
rect 3326 1584 3376 1618
rect 3326 1442 3370 1584
rect 3326 1406 3374 1442
rect 3326 1356 3376 1406
rect 3326 1318 3374 1356
rect 3410 1344 3420 1416
rect 3608 1344 3618 1416
rect 3326 1184 3370 1318
rect 3326 1176 3376 1184
rect 3658 1176 3898 1618
rect 3946 1340 3956 1420
rect 4138 1340 4148 1420
rect 3326 1140 4226 1176
rect 3326 1124 3376 1140
rect 3326 974 3370 1124
rect 3326 942 3374 974
rect 3658 972 3898 1140
rect 3656 942 3898 972
rect 3326 896 3898 942
rect 3326 882 3374 896
rect 3326 738 3370 882
rect 3656 878 3898 896
rect 3936 884 3946 958
rect 4148 884 4158 958
rect 3326 734 3376 738
rect 3658 734 3898 878
rect 3326 698 4232 734
rect 3326 678 3376 698
rect 3326 514 3370 678
rect 3326 488 3374 514
rect 3326 438 3376 488
rect 3326 428 3374 438
rect 3412 430 3422 502
rect 3610 430 3620 502
rect 3326 282 3370 428
rect 3424 426 3606 430
rect 3326 246 3376 282
rect 3658 246 3898 698
rect 5658 666 5692 828
rect 5732 822 5742 894
rect 5924 822 5934 894
rect 5972 820 6000 826
rect 5658 608 5966 666
rect 3944 426 3954 506
rect 4136 426 4146 506
rect 3326 210 4222 246
rect 3326 46 3370 210
rect 3326 28 3374 46
rect 3658 44 3898 210
rect 3656 28 3898 44
rect 5658 200 5692 608
rect 5728 434 5936 442
rect 5728 378 5738 434
rect 5928 378 5936 434
rect 5728 364 5936 378
rect 5972 200 6000 444
rect 5658 142 6000 200
rect 3326 -18 3898 28
rect 3326 -32 3374 -18
rect 3326 -200 3370 -32
rect 3656 -40 3898 -18
rect 3936 -32 3946 42
rect 4148 -32 4158 42
rect 3326 -206 3376 -200
rect 3658 -206 3898 -40
rect 3326 -242 4220 -206
rect 3326 -260 3376 -242
rect 3326 -402 3370 -260
rect 3658 -396 3898 -242
rect 3326 -582 3376 -402
rect 3424 -418 3606 -416
rect 3416 -478 3426 -418
rect 3608 -478 3618 -418
rect 3656 -458 3898 -396
rect 5658 -254 5692 142
rect 5730 -88 5740 -16
rect 5922 -88 5932 -16
rect 5972 -254 6000 142
rect 5658 -312 6000 -254
rect 3424 -486 3606 -478
rect 3656 -582 3706 -458
rect 3948 -488 3958 -418
rect 4138 -488 4148 -418
rect 5658 -480 5692 -312
rect 3954 -492 4140 -488
rect 5658 -544 5690 -480
rect 5658 -546 5698 -544
rect 3326 -650 3760 -582
rect 3962 -648 3972 -564
rect 4178 -648 4188 -564
rect 3534 -872 3634 -814
rect 3408 -970 3528 -902
rect 3408 -1382 3412 -970
rect 3502 -1382 3528 -970
rect 3408 -1404 3528 -1382
rect 3556 -1436 3612 -872
rect 3682 -902 3760 -650
rect 3920 -876 4022 -816
rect 3640 -1404 3760 -902
rect 3794 -980 3914 -904
rect 3788 -1378 3798 -980
rect 3882 -1378 3914 -980
rect 3794 -1404 3914 -1378
rect 3942 -1436 3998 -876
rect 4070 -904 4146 -648
rect 5658 -718 5692 -546
rect 5728 -564 5736 -462
rect 5928 -564 5936 -462
rect 5972 -718 6000 -312
rect 5658 -755 6000 -718
rect 4026 -1406 4146 -904
rect 4625 -776 6000 -755
rect 4625 -950 5692 -776
rect 1994 -1512 2224 -1496
rect 1994 -1874 2012 -1512
rect 2212 -1869 2224 -1512
rect 3534 -1712 3634 -1436
rect 3920 -1558 4020 -1436
rect 4343 -1540 4462 -1534
rect 3920 -1640 4343 -1558
rect 4343 -1665 4462 -1659
rect 3534 -1718 3982 -1712
rect 3534 -1822 3878 -1718
rect 3534 -1828 3982 -1822
rect 4625 -1869 4820 -950
rect 2212 -1874 4820 -1869
rect 1994 -2040 4820 -1874
rect 1996 -2041 4820 -2040
rect 5658 -1166 5692 -950
rect 5728 -996 5734 -944
rect 5930 -996 5936 -944
rect 5972 -1166 6000 -776
rect 6686 -842 6724 1756
rect 6758 1616 6768 1712
rect 6966 1616 6976 1712
rect 6760 1456 6770 1552
rect 6968 1456 6978 1552
rect 6764 1298 6774 1394
rect 6972 1298 6982 1394
rect 6762 1142 6772 1238
rect 6970 1142 6980 1238
rect 6764 982 6774 1078
rect 6972 982 6982 1078
rect 6762 826 6772 922
rect 6970 826 6980 922
rect 6764 666 6774 762
rect 6972 666 6982 762
rect 6762 510 6772 606
rect 6970 510 6980 606
rect 6760 350 6770 446
rect 6968 350 6978 446
rect 6762 194 6772 290
rect 6970 194 6980 290
rect 6762 34 6772 130
rect 6970 34 6980 130
rect 6762 -124 6772 -28
rect 6970 -124 6980 -28
rect 6764 -282 6774 -186
rect 6972 -282 6982 -186
rect 6762 -440 6772 -344
rect 6970 -440 6980 -344
rect 6764 -596 6774 -500
rect 6972 -596 6982 -500
rect 6762 -758 6772 -662
rect 6970 -758 6980 -662
rect 6762 -922 6772 -834
rect 6964 -922 6974 -834
rect 7014 -836 7052 2214
rect 7212 1926 7222 2392
rect 7610 2392 7988 2526
rect 7610 1926 7620 2392
rect 5658 -1224 6000 -1166
rect 5658 -1634 5692 -1224
rect 5728 -1398 5936 -1392
rect 5728 -1462 5736 -1398
rect 5928 -1462 5936 -1398
rect 5728 -1470 5936 -1462
rect 5972 -1634 6000 -1224
rect 5658 -1692 6000 -1634
rect 1996 -2042 4734 -2041
rect 2272 -2180 2422 -2042
rect 5658 -2088 5692 -1692
rect 5728 -1914 5734 -1860
rect 5928 -1914 5936 -1860
rect 5972 -2088 6000 -1692
rect 5658 -2146 6000 -2088
rect 2272 -2244 3818 -2180
rect 2326 -2254 3818 -2244
rect 2118 -2492 2128 -2292
rect 2180 -2492 2190 -2292
rect 2346 -2548 2422 -2254
rect 2578 -2492 2588 -2292
rect 2644 -2492 2654 -2292
rect 2808 -2546 2884 -2254
rect 3034 -2492 3044 -2292
rect 3100 -2492 3110 -2292
rect 3256 -2548 3332 -2254
rect 3492 -2492 3502 -2292
rect 3558 -2492 3568 -2292
rect 3724 -2548 3800 -2254
rect 3952 -2492 3962 -2292
rect 4018 -2492 4028 -2292
rect 5658 -2302 5692 -2146
rect 5728 -2314 5936 -2306
rect 5728 -2366 5738 -2314
rect 5928 -2366 5936 -2314
rect 5972 -2320 6000 -2146
rect 5728 -2374 5936 -2366
rect 5732 -2454 5932 -2374
rect 4126 -2516 7988 -2454
rect 4126 -2690 5128 -2516
rect 1988 -2702 5128 -2690
rect 1988 -2818 2132 -2702
rect 4010 -2736 5128 -2702
rect 7906 -2736 7988 -2516
rect 7908 -2814 7988 -2736
rect 1988 -3040 2228 -2818
rect 7908 -3040 7984 -2814
rect 1988 -3100 7984 -3040
<< via1 >>
rect 7222 2526 7610 2796
rect 3420 2272 3608 2344
rect 3956 2274 4138 2354
rect 6772 2246 6970 2342
rect 6772 2090 6970 2186
rect 6770 1930 6968 2026
rect 3946 1796 4148 1870
rect 6528 1788 6666 1876
rect 6770 1774 6968 1870
rect 3420 1344 3608 1416
rect 3956 1340 4138 1420
rect 3946 884 4148 958
rect 3422 430 3610 502
rect 5742 822 5924 894
rect 3954 426 4136 506
rect 5738 378 5928 434
rect 3946 -32 4148 42
rect 3426 -478 3608 -418
rect 5740 -88 5922 -16
rect 3958 -488 4138 -418
rect 3972 -648 4178 -564
rect 3412 -1382 3502 -970
rect 3798 -1378 3882 -980
rect 5736 -564 5928 -462
rect 2012 -1874 2212 -1512
rect 4343 -1659 4462 -1540
rect 3878 -1822 3982 -1718
rect 5734 -996 5930 -944
rect 6768 1616 6966 1712
rect 6770 1456 6968 1552
rect 6774 1298 6972 1394
rect 6772 1142 6970 1238
rect 6774 982 6972 1078
rect 6772 826 6970 922
rect 6774 666 6972 762
rect 6772 510 6970 606
rect 6770 350 6968 446
rect 6772 194 6970 290
rect 6772 34 6970 130
rect 6772 -124 6970 -28
rect 6774 -282 6972 -186
rect 6772 -440 6970 -344
rect 6774 -596 6972 -500
rect 6772 -758 6970 -662
rect 6772 -922 6964 -834
rect 7222 1926 7610 2526
rect 5736 -1462 5928 -1398
rect 5734 -1914 5928 -1860
rect 2128 -2492 2180 -2292
rect 2588 -2492 2644 -2292
rect 3044 -2492 3100 -2292
rect 3502 -2492 3558 -2292
rect 3962 -2492 4018 -2292
rect 5738 -2366 5928 -2314
rect 2132 -2736 4010 -2702
rect 2132 -2818 2228 -2736
rect 2228 -2818 4010 -2736
<< metal2 >>
rect 7222 2796 7610 2806
rect 3956 2354 4138 2364
rect 3420 2344 3608 2354
rect 3420 2262 3608 2272
rect 3956 2264 4138 2274
rect 6772 2342 6970 2352
rect 6772 2236 6970 2246
rect 6772 2186 7222 2198
rect 6970 2090 7222 2186
rect 6772 2082 7222 2090
rect 6772 2080 6970 2082
rect 6770 2026 6968 2036
rect 6770 1920 6968 1930
rect 7222 1916 7610 1926
rect 3946 1875 4148 1880
rect 6528 1876 6666 1886
rect 7226 1880 7430 1916
rect 3946 1870 6528 1875
rect 4148 1796 6528 1870
rect 3946 1789 6528 1796
rect 3946 1786 4148 1789
rect 3420 1416 3608 1426
rect 3420 1334 3608 1344
rect 3956 1420 4138 1430
rect 3956 1330 4138 1340
rect 3946 961 4148 968
rect 4305 961 4391 1789
rect 6666 1789 6721 1875
rect 6770 1870 7430 1880
rect 6528 1778 6666 1788
rect 6968 1774 7430 1870
rect 6770 1764 7430 1774
rect 6768 1712 6966 1722
rect 6768 1606 6966 1616
rect 7226 1562 7430 1764
rect 6770 1552 7430 1562
rect 6968 1456 7430 1552
rect 6770 1446 7430 1456
rect 6774 1394 6972 1404
rect 6774 1288 6972 1298
rect 7226 1248 7430 1446
rect 6772 1238 7430 1248
rect 6970 1142 7430 1238
rect 6772 1132 7430 1142
rect 6774 1078 6972 1088
rect 6774 972 6972 982
rect 3946 958 4391 961
rect 4148 884 4391 958
rect 7226 932 7430 1132
rect 6026 928 6198 930
rect 5744 904 6198 928
rect 3946 875 4391 884
rect 3946 874 4148 875
rect 3422 502 3610 512
rect 3422 420 3610 430
rect 3954 506 4136 516
rect 3954 416 4136 426
rect 3946 43 4148 52
rect 4305 43 4391 875
rect 5742 894 6198 904
rect 5924 822 6198 894
rect 5742 812 6198 822
rect 6772 922 7430 932
rect 6970 826 7430 922
rect 6772 820 7430 826
rect 6772 816 6970 820
rect 5744 782 6198 812
rect 5738 434 5928 444
rect 5738 368 5928 378
rect 3943 42 4391 43
rect 3943 -32 3946 42
rect 4148 -32 4391 42
rect 6026 18 6198 782
rect 6774 762 6972 772
rect 6774 656 6972 666
rect 6772 613 6970 616
rect 7226 613 7430 820
rect 6772 606 7430 613
rect 6970 510 7430 606
rect 6772 501 7430 510
rect 6772 500 6970 501
rect 6770 446 6968 456
rect 6770 340 6968 350
rect 6772 299 6970 300
rect 7226 299 7430 501
rect 6772 290 7430 299
rect 6970 194 7430 290
rect 6772 188 7430 194
rect 6772 184 6970 188
rect 6772 130 6970 140
rect 6772 24 6970 34
rect 3943 -43 4391 -32
rect 3426 -418 3608 -408
rect 3426 -488 3608 -478
rect 3958 -418 4138 -408
rect 3958 -498 4138 -488
rect 3972 -564 4178 -554
rect 4305 -564 4391 -43
rect 5740 -16 6198 18
rect 5922 -88 6198 -16
rect 5740 -128 6198 -88
rect 3970 -648 3972 -564
rect 4178 -648 4391 -564
rect 5736 -462 5928 -452
rect 5736 -574 5928 -564
rect 3970 -650 4391 -648
rect 3972 -658 4178 -650
rect 6026 -888 6198 -128
rect 6772 -21 6970 -18
rect 7226 -21 7430 188
rect 6772 -28 7430 -21
rect 6970 -124 7430 -28
rect 6772 -132 7430 -124
rect 6772 -134 6970 -132
rect 6774 -186 6972 -176
rect 6774 -292 6972 -282
rect 7226 -334 7430 -132
rect 6772 -344 7430 -334
rect 6970 -440 7430 -344
rect 6772 -450 7430 -440
rect 6774 -500 6972 -490
rect 6774 -606 6972 -596
rect 7226 -652 7430 -450
rect 6772 -662 7430 -652
rect 6970 -758 7430 -662
rect 6772 -764 7430 -758
rect 6772 -768 7358 -764
rect 6772 -824 6960 -816
rect 6772 -826 6964 -824
rect 5726 -944 6198 -888
rect 6766 -936 6772 -832
rect 6960 -832 6964 -826
rect 6960 -834 6970 -832
rect 6964 -922 6970 -834
rect 2926 -970 3898 -964
rect 2926 -1382 3412 -970
rect 3502 -980 3898 -970
rect 3502 -1378 3798 -980
rect 3882 -1378 3898 -980
rect 5726 -996 5734 -944
rect 5930 -996 6198 -944
rect 5726 -1034 6198 -996
rect 6026 -1216 6198 -1034
rect 6770 -940 6772 -936
rect 6960 -940 6970 -922
rect 6770 -1216 6970 -940
rect 3502 -1382 3898 -1378
rect 2926 -1394 3898 -1382
rect 2012 -1512 2212 -1502
rect 2926 -1834 3195 -1394
rect 3704 -1396 3898 -1394
rect 5736 -1388 5928 -1378
rect 5736 -1482 5928 -1472
rect 6026 -1468 7974 -1216
rect 4337 -1659 4343 -1540
rect 4462 -1543 4468 -1540
rect 4462 -1657 5005 -1543
rect 4462 -1659 4468 -1657
rect 3872 -1822 3878 -1718
rect 3982 -1726 4078 -1718
rect 4260 -1726 4476 -1718
rect 3982 -1822 4476 -1726
rect 2926 -1868 3194 -1834
rect 2012 -1884 2212 -1874
rect 2588 -2028 3558 -1868
rect 4372 -2012 4476 -1822
rect 4891 -1968 5005 -1657
rect 6026 -1816 6198 -1468
rect 5732 -1860 6198 -1816
rect 5732 -1914 5734 -1860
rect 5928 -1914 6198 -1860
rect 5732 -1962 6198 -1914
rect 2128 -2292 2180 -2282
rect 2128 -2586 2180 -2492
rect 2588 -2292 2644 -2028
rect 2588 -2502 2644 -2492
rect 3044 -2292 3100 -2282
rect 3044 -2502 3100 -2492
rect 3502 -2292 3558 -2028
rect 3502 -2502 3558 -2492
rect 3962 -2292 4018 -2282
rect 3962 -2502 4018 -2492
rect 3046 -2586 3098 -2502
rect 3964 -2586 4016 -2502
rect 2128 -2702 4016 -2586
rect 2128 -2818 2132 -2702
rect 4010 -2818 4016 -2702
rect 2132 -2828 4010 -2818
rect 4324 -3070 4524 -2012
rect 4848 -2882 5048 -1968
rect 5738 -2308 5928 -2298
rect 5738 -2386 5928 -2376
rect 4846 -3082 5048 -2882
<< via2 >>
rect 3420 2272 3608 2344
rect 3956 2274 4138 2354
rect 6772 2246 6970 2342
rect 6770 1930 6968 2026
rect 3420 1344 3608 1416
rect 3956 1340 4138 1420
rect 6768 1616 6966 1712
rect 6774 1298 6972 1394
rect 6774 982 6972 1078
rect 3422 430 3610 502
rect 3954 426 4136 506
rect 5738 378 5928 434
rect 6774 666 6972 762
rect 6770 350 6968 446
rect 6772 34 6970 130
rect 3426 -478 3608 -418
rect 3958 -488 4138 -418
rect 5736 -564 5928 -462
rect 6774 -282 6972 -186
rect 6774 -596 6972 -500
rect 6772 -834 6960 -826
rect 6772 -922 6960 -834
rect 6772 -940 6960 -922
rect 5736 -1398 5928 -1388
rect 5736 -1462 5928 -1398
rect 5736 -1472 5928 -1462
rect 5738 -2314 5928 -2308
rect 5738 -2366 5928 -2314
rect 5738 -2376 5928 -2366
<< metal3 >>
rect 3424 2349 3612 2384
rect 3956 2359 4136 2466
rect 3946 2354 4148 2359
rect 3410 2344 3618 2349
rect 3410 2272 3420 2344
rect 3608 2272 3618 2344
rect 3410 2267 3618 2272
rect 3946 2274 3956 2354
rect 4138 2274 4148 2354
rect 6772 2347 6974 2348
rect 3946 2269 4148 2274
rect 6762 2342 6980 2347
rect 3424 1421 3612 2267
rect 3956 1425 4136 2269
rect 6762 2246 6772 2342
rect 6970 2246 6980 2342
rect 6762 2241 6980 2246
rect 6772 2031 6974 2241
rect 6760 2026 6978 2031
rect 6760 1930 6770 2026
rect 6968 1930 6978 2026
rect 6760 1925 6978 1930
rect 6772 1717 6974 1925
rect 6758 1712 6976 1717
rect 6758 1616 6768 1712
rect 6966 1616 6976 1712
rect 6758 1611 6976 1616
rect 3410 1416 3618 1421
rect 3410 1344 3420 1416
rect 3608 1344 3618 1416
rect 3410 1339 3618 1344
rect 3946 1420 4148 1425
rect 3946 1340 3956 1420
rect 4138 1340 4148 1420
rect 6772 1399 6974 1611
rect 3424 507 3612 1339
rect 3946 1335 4148 1340
rect 6764 1394 6982 1399
rect 3956 511 4136 1335
rect 6764 1298 6774 1394
rect 6972 1298 6982 1394
rect 6764 1293 6982 1298
rect 6772 1083 6974 1293
rect 6764 1078 6982 1083
rect 6764 982 6774 1078
rect 6972 982 6982 1078
rect 6764 977 6982 982
rect 6772 767 6974 977
rect 6764 762 6982 767
rect 6764 666 6774 762
rect 6972 666 6982 762
rect 6764 661 6982 666
rect 3412 502 3620 507
rect 3412 430 3422 502
rect 3610 430 3620 502
rect 3412 425 3620 430
rect 3944 506 4146 511
rect 3944 426 3954 506
rect 4136 426 4146 506
rect 3424 -413 3612 425
rect 3944 421 4146 426
rect 5720 434 5944 472
rect 6772 451 6974 661
rect 3956 -413 4136 421
rect 5720 378 5738 434
rect 5928 378 5944 434
rect 3416 -418 3618 -413
rect 3416 -478 3426 -418
rect 3608 -478 3618 -418
rect 3416 -483 3618 -478
rect 3948 -418 4148 -413
rect 3948 -488 3958 -418
rect 4138 -488 4148 -418
rect 3948 -493 4148 -488
rect 5720 -462 5944 378
rect 6760 446 6978 451
rect 6760 350 6770 446
rect 6968 350 6978 446
rect 6760 345 6978 350
rect 6772 135 6974 345
rect 6762 130 6980 135
rect 6762 34 6772 130
rect 6970 34 6980 130
rect 6762 29 6980 34
rect 6772 -181 6974 29
rect 6764 -186 6982 -181
rect 6764 -282 6774 -186
rect 6972 -282 6982 -186
rect 6764 -287 6982 -282
rect 3956 -498 4136 -493
rect 5720 -564 5736 -462
rect 5928 -564 5944 -462
rect 6772 -495 6974 -287
rect 5720 -1388 5944 -564
rect 6764 -500 6982 -495
rect 6764 -596 6774 -500
rect 6972 -596 6982 -500
rect 6764 -601 6982 -596
rect 6772 -821 6974 -601
rect 6762 -826 6974 -821
rect 6762 -940 6772 -826
rect 6960 -922 6974 -826
rect 6960 -940 6970 -922
rect 6762 -945 6970 -940
rect 5720 -1472 5736 -1388
rect 5928 -1472 5944 -1388
rect 5720 -2308 5944 -1472
rect 5720 -2376 5738 -2308
rect 5928 -2376 5944 -2308
rect 5720 -2432 5944 -2376
use sky130_fd_pr__nfet_01v8_lvt_8TELWR  XM1
timestamp 1713292280
transform -1 0 3970 0 -1 -1154
box -246 -460 246 460
use sky130_fd_pr__nfet_01v8_lvt_8TELWR  XM2
timestamp 1713292280
transform -1 0 3584 0 -1 -1154
box -246 -460 246 460
use sky130_fd_pr__nfet_01v8_VWWVRL  XM3
timestamp 1713420874
transform -1 0 3073 0 -1 -2392
box -1083 -310 1083 310
use sky130_fd_pr__pfet_01v8_lvt_GW6ZVV  XM4
timestamp 1713292280
transform 0 1 3515 -1 0 921
box -1541 -319 1541 319
use sky130_fd_pr__pfet_01v8_lvt_GW6ZVV  XM5
timestamp 1713292280
transform 0 1 4047 -1 0 921
box -1541 -319 1541 319
use sky130_fd_pr__nfet_01v8_WWWVRA  XM7
timestamp 1713292280
transform 0 1 5832 -1 0 -742
box -1770 -310 1770 310
use sky130_fd_pr__pfet_01v8_lvt_ER3WAW  XM8
timestamp 1713292280
transform 0 1 6869 1 0 713
box -1747 -319 1747 319
<< labels >>
flabel metal1 1996 -3088 2196 -2888 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 1998 2690 2198 2890 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal2 2012 -1712 2212 -1512 0 FreeSans 256 0 0 0 VBIAS
port 0 nsew
flabel metal2 4324 -3070 4524 -2870 0 FreeSans 256 0 0 0 MINUS
port 2 nsew
flabel metal2 4846 -3082 5046 -2882 0 FreeSans 256 0 0 0 PLUS
port 3 nsew
flabel locali 2926 -2028 3195 -964 0 FreeSans 400 0 0 0 VX
flabel metal1 3496 -650 3760 -582 0 FreeSans 400 0 0 0 V2
flabel via1 4006 -642 4146 -580 0 FreeSans 400 0 0 0 V1
flabel metal2 7772 -1440 7972 -1240 0 FreeSans 256 0 0 0 VOUT
port 4 nsew
<< end >>
