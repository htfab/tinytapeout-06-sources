magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -1199 -1337 1199 1337
<< nmos >>
rect -1003 727 -803 1127
rect -745 727 -545 1127
rect -487 727 -287 1127
rect -229 727 -29 1127
rect 29 727 229 1127
rect 287 727 487 1127
rect 545 727 745 1127
rect 803 727 1003 1127
rect -1003 109 -803 509
rect -745 109 -545 509
rect -487 109 -287 509
rect -229 109 -29 509
rect 29 109 229 509
rect 287 109 487 509
rect 545 109 745 509
rect 803 109 1003 509
rect -1003 -509 -803 -109
rect -745 -509 -545 -109
rect -487 -509 -287 -109
rect -229 -509 -29 -109
rect 29 -509 229 -109
rect 287 -509 487 -109
rect 545 -509 745 -109
rect 803 -509 1003 -109
rect -1003 -1127 -803 -727
rect -745 -1127 -545 -727
rect -487 -1127 -287 -727
rect -229 -1127 -29 -727
rect 29 -1127 229 -727
rect 287 -1127 487 -727
rect 545 -1127 745 -727
rect 803 -1127 1003 -727
<< ndiff >>
rect -1061 1115 -1003 1127
rect -1061 739 -1049 1115
rect -1015 739 -1003 1115
rect -1061 727 -1003 739
rect -803 1115 -745 1127
rect -803 739 -791 1115
rect -757 739 -745 1115
rect -803 727 -745 739
rect -545 1115 -487 1127
rect -545 739 -533 1115
rect -499 739 -487 1115
rect -545 727 -487 739
rect -287 1115 -229 1127
rect -287 739 -275 1115
rect -241 739 -229 1115
rect -287 727 -229 739
rect -29 1115 29 1127
rect -29 739 -17 1115
rect 17 739 29 1115
rect -29 727 29 739
rect 229 1115 287 1127
rect 229 739 241 1115
rect 275 739 287 1115
rect 229 727 287 739
rect 487 1115 545 1127
rect 487 739 499 1115
rect 533 739 545 1115
rect 487 727 545 739
rect 745 1115 803 1127
rect 745 739 757 1115
rect 791 739 803 1115
rect 745 727 803 739
rect 1003 1115 1061 1127
rect 1003 739 1015 1115
rect 1049 739 1061 1115
rect 1003 727 1061 739
rect -1061 497 -1003 509
rect -1061 121 -1049 497
rect -1015 121 -1003 497
rect -1061 109 -1003 121
rect -803 497 -745 509
rect -803 121 -791 497
rect -757 121 -745 497
rect -803 109 -745 121
rect -545 497 -487 509
rect -545 121 -533 497
rect -499 121 -487 497
rect -545 109 -487 121
rect -287 497 -229 509
rect -287 121 -275 497
rect -241 121 -229 497
rect -287 109 -229 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 229 497 287 509
rect 229 121 241 497
rect 275 121 287 497
rect 229 109 287 121
rect 487 497 545 509
rect 487 121 499 497
rect 533 121 545 497
rect 487 109 545 121
rect 745 497 803 509
rect 745 121 757 497
rect 791 121 803 497
rect 745 109 803 121
rect 1003 497 1061 509
rect 1003 121 1015 497
rect 1049 121 1061 497
rect 1003 109 1061 121
rect -1061 -121 -1003 -109
rect -1061 -497 -1049 -121
rect -1015 -497 -1003 -121
rect -1061 -509 -1003 -497
rect -803 -121 -745 -109
rect -803 -497 -791 -121
rect -757 -497 -745 -121
rect -803 -509 -745 -497
rect -545 -121 -487 -109
rect -545 -497 -533 -121
rect -499 -497 -487 -121
rect -545 -509 -487 -497
rect -287 -121 -229 -109
rect -287 -497 -275 -121
rect -241 -497 -229 -121
rect -287 -509 -229 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 229 -121 287 -109
rect 229 -497 241 -121
rect 275 -497 287 -121
rect 229 -509 287 -497
rect 487 -121 545 -109
rect 487 -497 499 -121
rect 533 -497 545 -121
rect 487 -509 545 -497
rect 745 -121 803 -109
rect 745 -497 757 -121
rect 791 -497 803 -121
rect 745 -509 803 -497
rect 1003 -121 1061 -109
rect 1003 -497 1015 -121
rect 1049 -497 1061 -121
rect 1003 -509 1061 -497
rect -1061 -739 -1003 -727
rect -1061 -1115 -1049 -739
rect -1015 -1115 -1003 -739
rect -1061 -1127 -1003 -1115
rect -803 -739 -745 -727
rect -803 -1115 -791 -739
rect -757 -1115 -745 -739
rect -803 -1127 -745 -1115
rect -545 -739 -487 -727
rect -545 -1115 -533 -739
rect -499 -1115 -487 -739
rect -545 -1127 -487 -1115
rect -287 -739 -229 -727
rect -287 -1115 -275 -739
rect -241 -1115 -229 -739
rect -287 -1127 -229 -1115
rect -29 -739 29 -727
rect -29 -1115 -17 -739
rect 17 -1115 29 -739
rect -29 -1127 29 -1115
rect 229 -739 287 -727
rect 229 -1115 241 -739
rect 275 -1115 287 -739
rect 229 -1127 287 -1115
rect 487 -739 545 -727
rect 487 -1115 499 -739
rect 533 -1115 545 -739
rect 487 -1127 545 -1115
rect 745 -739 803 -727
rect 745 -1115 757 -739
rect 791 -1115 803 -739
rect 745 -1127 803 -1115
rect 1003 -739 1061 -727
rect 1003 -1115 1015 -739
rect 1049 -1115 1061 -739
rect 1003 -1127 1061 -1115
<< ndiffc >>
rect -1049 739 -1015 1115
rect -791 739 -757 1115
rect -533 739 -499 1115
rect -275 739 -241 1115
rect -17 739 17 1115
rect 241 739 275 1115
rect 499 739 533 1115
rect 757 739 791 1115
rect 1015 739 1049 1115
rect -1049 121 -1015 497
rect -791 121 -757 497
rect -533 121 -499 497
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect 499 121 533 497
rect 757 121 791 497
rect 1015 121 1049 497
rect -1049 -497 -1015 -121
rect -791 -497 -757 -121
rect -533 -497 -499 -121
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
rect 499 -497 533 -121
rect 757 -497 791 -121
rect 1015 -497 1049 -121
rect -1049 -1115 -1015 -739
rect -791 -1115 -757 -739
rect -533 -1115 -499 -739
rect -275 -1115 -241 -739
rect -17 -1115 17 -739
rect 241 -1115 275 -739
rect 499 -1115 533 -739
rect 757 -1115 791 -739
rect 1015 -1115 1049 -739
<< psubdiff >>
rect -1163 1267 1163 1301
rect -1163 1205 -1129 1267
rect 1129 1205 1163 1267
rect -1163 -1267 -1129 -1205
rect 1129 -1267 1163 -1205
rect -1163 -1301 -1067 -1267
rect 1067 -1301 1163 -1267
<< psubdiffcont >>
rect -1163 -1205 -1129 1205
rect 1129 -1205 1163 1205
rect -1067 -1301 1067 -1267
<< poly >>
rect -1003 1199 -803 1215
rect -1003 1165 -987 1199
rect -819 1165 -803 1199
rect -1003 1127 -803 1165
rect -745 1199 -545 1215
rect -745 1165 -729 1199
rect -561 1165 -545 1199
rect -745 1127 -545 1165
rect -487 1199 -287 1215
rect -487 1165 -471 1199
rect -303 1165 -287 1199
rect -487 1127 -287 1165
rect -229 1199 -29 1215
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect -229 1127 -29 1165
rect 29 1199 229 1215
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 29 1127 229 1165
rect 287 1199 487 1215
rect 287 1165 303 1199
rect 471 1165 487 1199
rect 287 1127 487 1165
rect 545 1199 745 1215
rect 545 1165 561 1199
rect 729 1165 745 1199
rect 545 1127 745 1165
rect 803 1199 1003 1215
rect 803 1165 819 1199
rect 987 1165 1003 1199
rect 803 1127 1003 1165
rect -1003 689 -803 727
rect -1003 655 -987 689
rect -819 655 -803 689
rect -1003 639 -803 655
rect -745 689 -545 727
rect -745 655 -729 689
rect -561 655 -545 689
rect -745 639 -545 655
rect -487 689 -287 727
rect -487 655 -471 689
rect -303 655 -287 689
rect -487 639 -287 655
rect -229 689 -29 727
rect -229 655 -213 689
rect -45 655 -29 689
rect -229 639 -29 655
rect 29 689 229 727
rect 29 655 45 689
rect 213 655 229 689
rect 29 639 229 655
rect 287 689 487 727
rect 287 655 303 689
rect 471 655 487 689
rect 287 639 487 655
rect 545 689 745 727
rect 545 655 561 689
rect 729 655 745 689
rect 545 639 745 655
rect 803 689 1003 727
rect 803 655 819 689
rect 987 655 1003 689
rect 803 639 1003 655
rect -1003 581 -803 597
rect -1003 547 -987 581
rect -819 547 -803 581
rect -1003 509 -803 547
rect -745 581 -545 597
rect -745 547 -729 581
rect -561 547 -545 581
rect -745 509 -545 547
rect -487 581 -287 597
rect -487 547 -471 581
rect -303 547 -287 581
rect -487 509 -287 547
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 509 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 509 229 547
rect 287 581 487 597
rect 287 547 303 581
rect 471 547 487 581
rect 287 509 487 547
rect 545 581 745 597
rect 545 547 561 581
rect 729 547 745 581
rect 545 509 745 547
rect 803 581 1003 597
rect 803 547 819 581
rect 987 547 1003 581
rect 803 509 1003 547
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect -1003 -547 -803 -509
rect -1003 -581 -987 -547
rect -819 -581 -803 -547
rect -1003 -597 -803 -581
rect -745 -547 -545 -509
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -745 -597 -545 -581
rect -487 -547 -287 -509
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -487 -597 -287 -581
rect -229 -547 -29 -509
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -509
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
rect 287 -547 487 -509
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 287 -597 487 -581
rect 545 -547 745 -509
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 545 -597 745 -581
rect 803 -547 1003 -509
rect 803 -581 819 -547
rect 987 -581 1003 -547
rect 803 -597 1003 -581
rect -1003 -655 -803 -639
rect -1003 -689 -987 -655
rect -819 -689 -803 -655
rect -1003 -727 -803 -689
rect -745 -655 -545 -639
rect -745 -689 -729 -655
rect -561 -689 -545 -655
rect -745 -727 -545 -689
rect -487 -655 -287 -639
rect -487 -689 -471 -655
rect -303 -689 -287 -655
rect -487 -727 -287 -689
rect -229 -655 -29 -639
rect -229 -689 -213 -655
rect -45 -689 -29 -655
rect -229 -727 -29 -689
rect 29 -655 229 -639
rect 29 -689 45 -655
rect 213 -689 229 -655
rect 29 -727 229 -689
rect 287 -655 487 -639
rect 287 -689 303 -655
rect 471 -689 487 -655
rect 287 -727 487 -689
rect 545 -655 745 -639
rect 545 -689 561 -655
rect 729 -689 745 -655
rect 545 -727 745 -689
rect 803 -655 1003 -639
rect 803 -689 819 -655
rect 987 -689 1003 -655
rect 803 -727 1003 -689
rect -1003 -1165 -803 -1127
rect -1003 -1199 -987 -1165
rect -819 -1199 -803 -1165
rect -1003 -1215 -803 -1199
rect -745 -1165 -545 -1127
rect -745 -1199 -729 -1165
rect -561 -1199 -545 -1165
rect -745 -1215 -545 -1199
rect -487 -1165 -287 -1127
rect -487 -1199 -471 -1165
rect -303 -1199 -287 -1165
rect -487 -1215 -287 -1199
rect -229 -1165 -29 -1127
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect -229 -1215 -29 -1199
rect 29 -1165 229 -1127
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 29 -1215 229 -1199
rect 287 -1165 487 -1127
rect 287 -1199 303 -1165
rect 471 -1199 487 -1165
rect 287 -1215 487 -1199
rect 545 -1165 745 -1127
rect 545 -1199 561 -1165
rect 729 -1199 745 -1165
rect 545 -1215 745 -1199
rect 803 -1165 1003 -1127
rect 803 -1199 819 -1165
rect 987 -1199 1003 -1165
rect 803 -1215 1003 -1199
<< polycont >>
rect -987 1165 -819 1199
rect -729 1165 -561 1199
rect -471 1165 -303 1199
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect 303 1165 471 1199
rect 561 1165 729 1199
rect 819 1165 987 1199
rect -987 655 -819 689
rect -729 655 -561 689
rect -471 655 -303 689
rect -213 655 -45 689
rect 45 655 213 689
rect 303 655 471 689
rect 561 655 729 689
rect 819 655 987 689
rect -987 547 -819 581
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect 819 547 987 581
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect -987 -581 -819 -547
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
rect 819 -581 987 -547
rect -987 -689 -819 -655
rect -729 -689 -561 -655
rect -471 -689 -303 -655
rect -213 -689 -45 -655
rect 45 -689 213 -655
rect 303 -689 471 -655
rect 561 -689 729 -655
rect 819 -689 987 -655
rect -987 -1199 -819 -1165
rect -729 -1199 -561 -1165
rect -471 -1199 -303 -1165
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
rect 303 -1199 471 -1165
rect 561 -1199 729 -1165
rect 819 -1199 987 -1165
<< locali >>
rect -1163 1205 -1129 1301
rect 1129 1205 1163 1301
rect -1003 1165 -987 1199
rect -819 1165 -803 1199
rect -745 1165 -729 1199
rect -561 1165 -545 1199
rect -487 1165 -471 1199
rect -303 1165 -287 1199
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 287 1165 303 1199
rect 471 1165 487 1199
rect 545 1165 561 1199
rect 729 1165 745 1199
rect 803 1165 819 1199
rect 987 1165 1003 1199
rect -1049 1115 -1015 1131
rect -1049 723 -1015 739
rect -791 1115 -757 1131
rect -791 723 -757 739
rect -533 1115 -499 1131
rect -533 723 -499 739
rect -275 1115 -241 1131
rect -275 723 -241 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 241 1115 275 1131
rect 241 723 275 739
rect 499 1115 533 1131
rect 499 723 533 739
rect 757 1115 791 1131
rect 757 723 791 739
rect 1015 1115 1049 1131
rect 1015 723 1049 739
rect -1003 655 -987 689
rect -819 655 -803 689
rect -745 655 -729 689
rect -561 655 -545 689
rect -487 655 -471 689
rect -303 655 -287 689
rect -229 655 -213 689
rect -45 655 -29 689
rect 29 655 45 689
rect 213 655 229 689
rect 287 655 303 689
rect 471 655 487 689
rect 545 655 561 689
rect 729 655 745 689
rect 803 655 819 689
rect 987 655 1003 689
rect -1003 547 -987 581
rect -819 547 -803 581
rect -745 547 -729 581
rect -561 547 -545 581
rect -487 547 -471 581
rect -303 547 -287 581
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect 287 547 303 581
rect 471 547 487 581
rect 545 547 561 581
rect 729 547 745 581
rect 803 547 819 581
rect 987 547 1003 581
rect -1049 497 -1015 513
rect -1049 105 -1015 121
rect -791 497 -757 513
rect -791 105 -757 121
rect -533 497 -499 513
rect -533 105 -499 121
rect -275 497 -241 513
rect -275 105 -241 121
rect -17 497 17 513
rect -17 105 17 121
rect 241 497 275 513
rect 241 105 275 121
rect 499 497 533 513
rect 499 105 533 121
rect 757 497 791 513
rect 757 105 791 121
rect 1015 497 1049 513
rect 1015 105 1049 121
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect -1049 -121 -1015 -105
rect -1049 -513 -1015 -497
rect -791 -121 -757 -105
rect -791 -513 -757 -497
rect -533 -121 -499 -105
rect -533 -513 -499 -497
rect -275 -121 -241 -105
rect -275 -513 -241 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 241 -121 275 -105
rect 241 -513 275 -497
rect 499 -121 533 -105
rect 499 -513 533 -497
rect 757 -121 791 -105
rect 757 -513 791 -497
rect 1015 -121 1049 -105
rect 1015 -513 1049 -497
rect -1003 -581 -987 -547
rect -819 -581 -803 -547
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 803 -581 819 -547
rect 987 -581 1003 -547
rect -1003 -689 -987 -655
rect -819 -689 -803 -655
rect -745 -689 -729 -655
rect -561 -689 -545 -655
rect -487 -689 -471 -655
rect -303 -689 -287 -655
rect -229 -689 -213 -655
rect -45 -689 -29 -655
rect 29 -689 45 -655
rect 213 -689 229 -655
rect 287 -689 303 -655
rect 471 -689 487 -655
rect 545 -689 561 -655
rect 729 -689 745 -655
rect 803 -689 819 -655
rect 987 -689 1003 -655
rect -1049 -739 -1015 -723
rect -1049 -1131 -1015 -1115
rect -791 -739 -757 -723
rect -791 -1131 -757 -1115
rect -533 -739 -499 -723
rect -533 -1131 -499 -1115
rect -275 -739 -241 -723
rect -275 -1131 -241 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 241 -739 275 -723
rect 241 -1131 275 -1115
rect 499 -739 533 -723
rect 499 -1131 533 -1115
rect 757 -739 791 -723
rect 757 -1131 791 -1115
rect 1015 -739 1049 -723
rect 1015 -1131 1049 -1115
rect -1003 -1199 -987 -1165
rect -819 -1199 -803 -1165
rect -745 -1199 -729 -1165
rect -561 -1199 -545 -1165
rect -487 -1199 -471 -1165
rect -303 -1199 -287 -1165
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 287 -1199 303 -1165
rect 471 -1199 487 -1165
rect 545 -1199 561 -1165
rect 729 -1199 745 -1165
rect 803 -1199 819 -1165
rect 987 -1199 1003 -1165
rect -1163 -1301 -1067 -1267
rect 1067 -1301 1163 -1267
<< viali >>
rect -1129 1267 1129 1301
rect -987 1165 -819 1199
rect -729 1165 -561 1199
rect -471 1165 -303 1199
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect 303 1165 471 1199
rect 561 1165 729 1199
rect 819 1165 987 1199
rect -1049 948 -1015 1098
rect -791 756 -757 906
rect -533 948 -499 1098
rect -275 756 -241 906
rect -17 948 17 1098
rect 241 756 275 906
rect 499 948 533 1098
rect 757 756 791 906
rect 1015 948 1049 1098
rect -987 655 -819 689
rect -729 655 -561 689
rect -471 655 -303 689
rect -213 655 -45 689
rect 45 655 213 689
rect 303 655 471 689
rect 561 655 729 689
rect 819 655 987 689
rect -987 547 -819 581
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect 819 547 987 581
rect -1049 330 -1015 480
rect -791 138 -757 288
rect -533 330 -499 480
rect -275 138 -241 288
rect -17 330 17 480
rect 241 138 275 288
rect 499 330 533 480
rect 757 138 791 288
rect 1015 330 1049 480
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect -1163 -1205 -1129 -253
rect -1049 -288 -1015 -138
rect -791 -480 -757 -330
rect -533 -288 -499 -138
rect -275 -480 -241 -330
rect -17 -288 17 -138
rect 241 -480 275 -330
rect 499 -288 533 -138
rect 757 -480 791 -330
rect 1015 -288 1049 -138
rect -987 -581 -819 -547
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
rect 819 -581 987 -547
rect -987 -689 -819 -655
rect -729 -689 -561 -655
rect -471 -689 -303 -655
rect -213 -689 -45 -655
rect 45 -689 213 -655
rect 303 -689 471 -655
rect 561 -689 729 -655
rect 819 -689 987 -655
rect -1049 -906 -1015 -756
rect -791 -1098 -757 -948
rect -533 -906 -499 -756
rect -275 -1098 -241 -948
rect -17 -906 17 -756
rect 241 -1098 275 -948
rect 499 -906 533 -756
rect 757 -1098 791 -948
rect 1015 -906 1049 -756
rect -987 -1199 -819 -1165
rect -729 -1199 -561 -1165
rect -471 -1199 -303 -1165
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
rect 303 -1199 471 -1165
rect 561 -1199 729 -1165
rect 819 -1199 987 -1165
rect -1163 -1267 -1129 -1205
rect 1129 -1205 1163 -253
rect 1129 -1267 1163 -1205
<< metal1 >>
rect -1141 1301 1141 1307
rect -1141 1267 -1129 1301
rect 1129 1267 1141 1301
rect -1141 1261 1141 1267
rect -999 1199 -807 1205
rect -999 1165 -987 1199
rect -819 1165 -807 1199
rect -999 1159 -807 1165
rect -741 1199 -549 1205
rect -741 1165 -729 1199
rect -561 1165 -549 1199
rect -741 1159 -549 1165
rect -483 1199 -291 1205
rect -483 1165 -471 1199
rect -303 1165 -291 1199
rect -483 1159 -291 1165
rect -225 1199 -33 1205
rect -225 1165 -213 1199
rect -45 1165 -33 1199
rect -225 1159 -33 1165
rect 33 1199 225 1205
rect 33 1165 45 1199
rect 213 1165 225 1199
rect 33 1159 225 1165
rect 291 1199 483 1205
rect 291 1165 303 1199
rect 471 1165 483 1199
rect 291 1159 483 1165
rect 549 1199 741 1205
rect 549 1165 561 1199
rect 729 1165 741 1199
rect 549 1159 741 1165
rect 807 1199 999 1205
rect 807 1165 819 1199
rect 987 1165 999 1199
rect 807 1159 999 1165
rect -1055 1098 -1009 1110
rect -1055 948 -1049 1098
rect -1015 948 -1009 1098
rect -1055 936 -1009 948
rect -539 1098 -493 1110
rect -539 948 -533 1098
rect -499 948 -493 1098
rect -539 936 -493 948
rect -23 1098 23 1110
rect -23 948 -17 1098
rect 17 948 23 1098
rect -23 936 23 948
rect 493 1098 539 1110
rect 493 948 499 1098
rect 533 948 539 1098
rect 493 936 539 948
rect 1009 1098 1055 1110
rect 1009 948 1015 1098
rect 1049 948 1055 1098
rect 1009 936 1055 948
rect -797 906 -751 918
rect -797 756 -791 906
rect -757 756 -751 906
rect -797 744 -751 756
rect -281 906 -235 918
rect -281 756 -275 906
rect -241 756 -235 906
rect -281 744 -235 756
rect 235 906 281 918
rect 235 756 241 906
rect 275 756 281 906
rect 235 744 281 756
rect 751 906 797 918
rect 751 756 757 906
rect 791 756 797 906
rect 751 744 797 756
rect -999 689 -807 695
rect -999 655 -987 689
rect -819 655 -807 689
rect -999 649 -807 655
rect -741 689 -549 695
rect -741 655 -729 689
rect -561 655 -549 689
rect -741 649 -549 655
rect -483 689 -291 695
rect -483 655 -471 689
rect -303 655 -291 689
rect -483 649 -291 655
rect -225 689 -33 695
rect -225 655 -213 689
rect -45 655 -33 689
rect -225 649 -33 655
rect 33 689 225 695
rect 33 655 45 689
rect 213 655 225 689
rect 33 649 225 655
rect 291 689 483 695
rect 291 655 303 689
rect 471 655 483 689
rect 291 649 483 655
rect 549 689 741 695
rect 549 655 561 689
rect 729 655 741 689
rect 549 649 741 655
rect 807 689 999 695
rect 807 655 819 689
rect 987 655 999 689
rect 807 649 999 655
rect -999 581 -807 587
rect -999 547 -987 581
rect -819 547 -807 581
rect -999 541 -807 547
rect -741 581 -549 587
rect -741 547 -729 581
rect -561 547 -549 581
rect -741 541 -549 547
rect -483 581 -291 587
rect -483 547 -471 581
rect -303 547 -291 581
rect -483 541 -291 547
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect 291 581 483 587
rect 291 547 303 581
rect 471 547 483 581
rect 291 541 483 547
rect 549 581 741 587
rect 549 547 561 581
rect 729 547 741 581
rect 549 541 741 547
rect 807 581 999 587
rect 807 547 819 581
rect 987 547 999 581
rect 807 541 999 547
rect -1055 480 -1009 492
rect -1055 330 -1049 480
rect -1015 330 -1009 480
rect -1055 318 -1009 330
rect -539 480 -493 492
rect -539 330 -533 480
rect -499 330 -493 480
rect -539 318 -493 330
rect -23 480 23 492
rect -23 330 -17 480
rect 17 330 23 480
rect -23 318 23 330
rect 493 480 539 492
rect 493 330 499 480
rect 533 330 539 480
rect 493 318 539 330
rect 1009 480 1055 492
rect 1009 330 1015 480
rect 1049 330 1055 480
rect 1009 318 1055 330
rect -797 288 -751 300
rect -797 138 -791 288
rect -757 138 -751 288
rect -797 126 -751 138
rect -281 288 -235 300
rect -281 138 -275 288
rect -241 138 -235 288
rect -281 126 -235 138
rect 235 288 281 300
rect 235 138 241 288
rect 275 138 281 288
rect 235 126 281 138
rect 751 288 797 300
rect 751 138 757 288
rect 791 138 797 288
rect 751 126 797 138
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect -1055 -138 -1009 -126
rect -1169 -253 -1123 -241
rect -1169 -1267 -1163 -253
rect -1129 -1267 -1123 -253
rect -1055 -288 -1049 -138
rect -1015 -288 -1009 -138
rect -1055 -300 -1009 -288
rect -539 -138 -493 -126
rect -539 -288 -533 -138
rect -499 -288 -493 -138
rect -539 -300 -493 -288
rect -23 -138 23 -126
rect -23 -288 -17 -138
rect 17 -288 23 -138
rect -23 -300 23 -288
rect 493 -138 539 -126
rect 493 -288 499 -138
rect 533 -288 539 -138
rect 493 -300 539 -288
rect 1009 -138 1055 -126
rect 1009 -288 1015 -138
rect 1049 -288 1055 -138
rect 1009 -300 1055 -288
rect 1123 -253 1169 -241
rect -797 -330 -751 -318
rect -797 -480 -791 -330
rect -757 -480 -751 -330
rect -797 -492 -751 -480
rect -281 -330 -235 -318
rect -281 -480 -275 -330
rect -241 -480 -235 -330
rect -281 -492 -235 -480
rect 235 -330 281 -318
rect 235 -480 241 -330
rect 275 -480 281 -330
rect 235 -492 281 -480
rect 751 -330 797 -318
rect 751 -480 757 -330
rect 791 -480 797 -330
rect 751 -492 797 -480
rect -999 -547 -807 -541
rect -999 -581 -987 -547
rect -819 -581 -807 -547
rect -999 -587 -807 -581
rect -741 -547 -549 -541
rect -741 -581 -729 -547
rect -561 -581 -549 -547
rect -741 -587 -549 -581
rect -483 -547 -291 -541
rect -483 -581 -471 -547
rect -303 -581 -291 -547
rect -483 -587 -291 -581
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
rect 291 -547 483 -541
rect 291 -581 303 -547
rect 471 -581 483 -547
rect 291 -587 483 -581
rect 549 -547 741 -541
rect 549 -581 561 -547
rect 729 -581 741 -547
rect 549 -587 741 -581
rect 807 -547 999 -541
rect 807 -581 819 -547
rect 987 -581 999 -547
rect 807 -587 999 -581
rect -999 -655 -807 -649
rect -999 -689 -987 -655
rect -819 -689 -807 -655
rect -999 -695 -807 -689
rect -741 -655 -549 -649
rect -741 -689 -729 -655
rect -561 -689 -549 -655
rect -741 -695 -549 -689
rect -483 -655 -291 -649
rect -483 -689 -471 -655
rect -303 -689 -291 -655
rect -483 -695 -291 -689
rect -225 -655 -33 -649
rect -225 -689 -213 -655
rect -45 -689 -33 -655
rect -225 -695 -33 -689
rect 33 -655 225 -649
rect 33 -689 45 -655
rect 213 -689 225 -655
rect 33 -695 225 -689
rect 291 -655 483 -649
rect 291 -689 303 -655
rect 471 -689 483 -655
rect 291 -695 483 -689
rect 549 -655 741 -649
rect 549 -689 561 -655
rect 729 -689 741 -655
rect 549 -695 741 -689
rect 807 -655 999 -649
rect 807 -689 819 -655
rect 987 -689 999 -655
rect 807 -695 999 -689
rect -1055 -756 -1009 -744
rect -1055 -906 -1049 -756
rect -1015 -906 -1009 -756
rect -1055 -918 -1009 -906
rect -539 -756 -493 -744
rect -539 -906 -533 -756
rect -499 -906 -493 -756
rect -539 -918 -493 -906
rect -23 -756 23 -744
rect -23 -906 -17 -756
rect 17 -906 23 -756
rect -23 -918 23 -906
rect 493 -756 539 -744
rect 493 -906 499 -756
rect 533 -906 539 -756
rect 493 -918 539 -906
rect 1009 -756 1055 -744
rect 1009 -906 1015 -756
rect 1049 -906 1055 -756
rect 1009 -918 1055 -906
rect -797 -948 -751 -936
rect -797 -1098 -791 -948
rect -757 -1098 -751 -948
rect -797 -1110 -751 -1098
rect -281 -948 -235 -936
rect -281 -1098 -275 -948
rect -241 -1098 -235 -948
rect -281 -1110 -235 -1098
rect 235 -948 281 -936
rect 235 -1098 241 -948
rect 275 -1098 281 -948
rect 235 -1110 281 -1098
rect 751 -948 797 -936
rect 751 -1098 757 -948
rect 791 -1098 797 -948
rect 751 -1110 797 -1098
rect -999 -1165 -807 -1159
rect -999 -1199 -987 -1165
rect -819 -1199 -807 -1165
rect -999 -1205 -807 -1199
rect -741 -1165 -549 -1159
rect -741 -1199 -729 -1165
rect -561 -1199 -549 -1165
rect -741 -1205 -549 -1199
rect -483 -1165 -291 -1159
rect -483 -1199 -471 -1165
rect -303 -1199 -291 -1165
rect -483 -1205 -291 -1199
rect -225 -1165 -33 -1159
rect -225 -1199 -213 -1165
rect -45 -1199 -33 -1165
rect -225 -1205 -33 -1199
rect 33 -1165 225 -1159
rect 33 -1199 45 -1165
rect 213 -1199 225 -1165
rect 33 -1205 225 -1199
rect 291 -1165 483 -1159
rect 291 -1199 303 -1165
rect 471 -1199 483 -1165
rect 291 -1205 483 -1199
rect 549 -1165 741 -1159
rect 549 -1199 561 -1165
rect 729 -1199 741 -1165
rect 549 -1205 741 -1199
rect 807 -1165 999 -1159
rect 807 -1199 819 -1165
rect 987 -1199 999 -1165
rect 807 -1205 999 -1199
rect -1169 -1279 -1123 -1267
rect 1123 -1267 1129 -253
rect 1163 -1267 1169 -253
rect 1123 -1279 1169 -1267
<< properties >>
string FIXED_BBOX -1146 -1284 1146 1284
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
