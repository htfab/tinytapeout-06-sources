** sch_path: /home/james/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-programmable-thing/xschem/inverter.sch
.subckt inverter VDD VSS OUT IN
*.PININFO VDD:B VSS:B IN:I OUT:O
XM1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=1
XM2 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=10 nf=1 m=1
.ends
.end
