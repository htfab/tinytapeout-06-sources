* NGSPICE file created from opamp_parax.ext - technology: sky130A

.subckt opamp_parax VBIAS VDD MINUS PLUS VOUT VSS
X0 VDD.t39 V1.t7 VOUT.t14 VDD.t38 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 VOUT.t24 VBIAS.t0 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X2 VDD.t37 V1.t8 VOUT.t12 VDD.t36 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 V1.t3 V2.t13 VDD.t48 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X4 VDD.t35 V1.t9 VOUT.t8 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 VOUT.t20 VBIAS.t1 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X6 VOUT.t13 V1.t10 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 VSS.t15 VBIAS.t2 VOUT.t22 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X8 VDD.t42 V2.t14 V1.t1 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X9 VDD.t44 V2.t11 V2.t12 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X10 V2.t10 V2.t9 VDD.t45 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X11 VSS.t14 VBIAS.t3 VOUT.t25 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X12 V2.t8 V2.t7 VDD.t46 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X13 VDD.t49 V2.t15 V1.t4 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X14 V1.t0 V2.t16 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X15 VDD.t51 V2.t5 V2.t6 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X16 V2.t0 MINUS.t0 a_2586_n2492# VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X17 VOUT.t26 VBIAS.t4 VSS.t12 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X18 VSS.t4 VBIAS.t5 VOUT.t23 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X19 VOUT.t9 V1.t11 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X20 V1.t6 PLUS.t0 a_2586_n2492# VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X21 VSS.t11 VBIAS.t6 a_2586_n2492# VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X22 V2.t4 V2.t3 VDD.t52 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X23 VOUT.t21 VBIAS.t7 VSS.t9 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X24 VDD.t29 V1.t12 VOUT.t15 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 VOUT.t10 V1.t13 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 VDD.t47 V2.t17 V1.t2 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X27 a_2586_n2492# VBIAS.t8 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X28 VDD.t25 V1.t14 VOUT.t11 VDD.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X29 VOUT.t3 V1.t15 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X30 VOUT.t2 V1.t16 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 VOUT.t16 V1.t17 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X32 VDD.t17 V1.t18 VOUT.t17 VDD.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X33 VDD.t15 V1.t19 VOUT.t0 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X34 VSS.t6 VBIAS.t9 a_2586_n2492# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X35 a_2586_n2492# VBIAS.t10 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X36 VOUT.t18 V1.t20 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X37 VDD.t11 V1.t21 VOUT.t1 VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 VOUT.t19 V1.t22 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X39 V1.t5 V2.t18 VDD.t53 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X40 VOUT.t4 V1.t23 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X41 VOUT.t7 V1.t24 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X42 VDD.t3 V1.t25 VOUT.t6 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 VDD.t50 V2.t1 V2.t2 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X44 VDD.t1 V1.t26 VOUT.t5 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
R0 V1.n7 V1.t18 240.815
R1 V1.n6 V1.t18 240.815
R2 V1.n4 V1.t9 240.351
R3 V1.t22 V1.n6 240.349
R4 V1.n7 V1.t22 240.349
R5 V1.t8 V1.n6 240.349
R6 V1.n7 V1.t8 240.349
R7 V1.n6 V1.t10 240.349
R8 V1.t10 V1.n7 240.349
R9 V1.n5 V1.t25 240.349
R10 V1.t25 V1.n7 240.349
R11 V1.t11 V1.n5 240.349
R12 V1.n8 V1.t11 240.349
R13 V1.t26 V1.n5 240.349
R14 V1.n8 V1.t26 240.349
R15 V1.n5 V1.t17 240.349
R16 V1.t17 V1.n8 240.349
R17 V1.n3 V1.t14 240.349
R18 V1.t14 V1.n8 240.349
R19 V1.t24 V1.n3 240.349
R20 V1.n9 V1.t24 240.349
R21 V1.t19 V1.n3 240.349
R22 V1.n9 V1.t19 240.349
R23 V1.n3 V1.t15 240.349
R24 V1.t15 V1.n9 240.349
R25 V1.n4 V1.t21 240.349
R26 V1.t21 V1.n9 240.349
R27 V1.t16 V1.n4 240.349
R28 V1.n0 V1.t16 240.349
R29 V1.t7 V1.n4 240.349
R30 V1.n0 V1.t7 240.349
R31 V1.n4 V1.t23 240.349
R32 V1.t23 V1.n0 240.349
R33 V1.n0 V1.t9 240.349
R34 V1.n1 V1.t12 119.487
R35 V1.n0 V1.t13 240.349
R36 V1.t13 V1.n4 240.353
R37 V1.n2 V1.n10 201.577
R38 V1.n2 V1.n11 201.576
R39 V1 V1.n12 201.575
R40 V1.n0 V1.t20 119.716
R41 V1 V1.t6 36.9223
R42 V1.n10 V1.t1 28.5655
R43 V1.n10 V1.t3 28.5655
R44 V1.n11 V1.t4 28.5655
R45 V1.n11 V1.t0 28.5655
R46 V1.n12 V1.t2 28.5655
R47 V1.n12 V1.t5 28.5655
R48 V1.n2 V1.n4 5.50039
R49 V1 V1.n2 3.54145
R50 V1.n8 V1.n7 2.80313
R51 V1.n4 V1.n1 3.66886
R52 V1.n1 V1.n0 2.77966
R53 V1.n0 V1.n9 1.86892
R54 V1.n9 V1.n8 1.86892
R55 V1.n5 V1.n6 1.86892
R56 V1.n3 V1.n5 1.86892
R57 V1.n4 V1.n3 1.86892
R58 VOUT.n1 VOUT.t18 231.496
R59 VOUT.n18 VOUT.t17 229.726
R60 VOUT.n5 VOUT.n4 202.861
R61 VOUT.n7 VOUT.n6 202.861
R62 VOUT.n9 VOUT.n8 202.861
R63 VOUT.n15 VOUT.n14 202.861
R64 VOUT.n17 VOUT.n16 202.861
R65 VOUT.n13 VOUT.n12 202.858
R66 VOUT.n3 VOUT.n2 202.857
R67 VOUT.n1 VOUT.n0 202.857
R68 VOUT.n11 VOUT.n10 202.857
R69 VOUT.n21 VOUT.t24 86.0456
R70 VOUT.n24 VOUT.n23 68.2924
R71 VOUT.n21 VOUT.n20 67.986
R72 VOUT.n22 VOUT.n19 67.9839
R73 VOUT.n0 VOUT.t15 28.5655
R74 VOUT.n0 VOUT.t10 28.5655
R75 VOUT.n2 VOUT.t8 28.5655
R76 VOUT.n2 VOUT.t4 28.5655
R77 VOUT.n4 VOUT.t14 28.5655
R78 VOUT.n4 VOUT.t2 28.5655
R79 VOUT.n6 VOUT.t1 28.5655
R80 VOUT.n6 VOUT.t3 28.5655
R81 VOUT.n8 VOUT.t0 28.5655
R82 VOUT.n8 VOUT.t7 28.5655
R83 VOUT.n10 VOUT.t11 28.5655
R84 VOUT.n10 VOUT.t16 28.5655
R85 VOUT.n12 VOUT.t5 28.5655
R86 VOUT.n12 VOUT.t9 28.5655
R87 VOUT.n14 VOUT.t6 28.5655
R88 VOUT.n14 VOUT.t13 28.5655
R89 VOUT.n16 VOUT.t12 28.5655
R90 VOUT.n16 VOUT.t19 28.5655
R91 VOUT.n23 VOUT.t23 17.4005
R92 VOUT.n23 VOUT.t21 17.4005
R93 VOUT.n19 VOUT.t22 17.4005
R94 VOUT.n19 VOUT.t26 17.4005
R95 VOUT.n20 VOUT.t25 17.4005
R96 VOUT.n20 VOUT.t20 17.4005
R97 VOUT.n18 VOUT.n17 1.78343
R98 VOUT.n22 VOUT.n21 0.65893
R99 VOUT VOUT.n25 0.447921
R100 VOUT.n25 VOUT.n24 0.376492
R101 VOUT.n25 VOUT.n18 0.208625
R102 VOUT.n24 VOUT.n22 0.18582
R103 VOUT.n5 VOUT.n3 0.0744901
R104 VOUT.n7 VOUT.n5 0.0740248
R105 VOUT.n9 VOUT.n7 0.0740248
R106 VOUT.n11 VOUT.n9 0.0740248
R107 VOUT.n13 VOUT.n11 0.0740248
R108 VOUT.n15 VOUT.n13 0.0740248
R109 VOUT.n3 VOUT.n1 0.0735594
R110 VOUT.n17 VOUT.n15 0.0735594
R111 VDD.n40 VDD.n36 6857.65
R112 VDD.n38 VDD.n36 6857.65
R113 VDD.n38 VDD.n35 6857.65
R114 VDD.n40 VDD.n35 6857.65
R115 VDD.n12 VDD.n9 6130.59
R116 VDD.n67 VDD.n8 6130.59
R117 VDD.n64 VDD.n63 5191.76
R118 VDD.n63 VDD.n10 5191.76
R119 VDD.n64 VDD.n9 938.823
R120 VDD.n65 VDD.n64 938.823
R121 VDD.n60 VDD.n10 938.823
R122 VDD.n10 VDD.n8 938.823
R123 VDD.n54 VDD.n11 553.788
R124 VDD.n58 VDD.n11 553.788
R125 VDD.n40 VDD.t12 318.216
R126 VDD.t16 VDD.n38 318.216
R127 VDD.t12 VDD.t28 235.267
R128 VDD.t28 VDD.t26 235.267
R129 VDD.t26 VDD.t34 235.267
R130 VDD.t34 VDD.t6 235.267
R131 VDD.t6 VDD.t38 235.267
R132 VDD.t38 VDD.t20 235.267
R133 VDD.t20 VDD.t10 235.267
R134 VDD.t10 VDD.t22 235.267
R135 VDD.t22 VDD.t14 235.267
R136 VDD.t4 VDD.t24 235.267
R137 VDD.t24 VDD.t18 235.267
R138 VDD.t18 VDD.t0 235.267
R139 VDD.t0 VDD.t30 235.267
R140 VDD.t30 VDD.t2 235.267
R141 VDD.t2 VDD.t32 235.267
R142 VDD.t32 VDD.t36 235.267
R143 VDD.t36 VDD.t8 235.267
R144 VDD.t8 VDD.t16 235.267
R145 VDD.n47 VDD.t53 231.662
R146 VDD.n1 VDD.t46 231.653
R147 VDD.n50 VDD.t42 228.226
R148 VDD.n4 VDD.t50 228.222
R149 VDD.n47 VDD.n46 202.858
R150 VDD.n1 VDD.n0 202.857
R151 VDD.n3 VDD.n2 202.857
R152 VDD.n49 VDD.n48 202.857
R153 VDD.n24 VDD.n23 201.73
R154 VDD.n25 VDD.n21 201.548
R155 VDD.n26 VDD.n20 201.548
R156 VDD.n27 VDD.n19 201.544
R157 VDD.n28 VDD.n18 201.544
R158 VDD.n31 VDD.n15 201.536
R159 VDD.n30 VDD.n16 201.536
R160 VDD.n24 VDD.n22 201.536
R161 VDD.n29 VDD.n17 201.535
R162 VDD.n32 VDD.n14 201.529
R163 VDD.t14 VDD.n39 117.633
R164 VDD.n39 VDD.t4 117.633
R165 VDD.n37 VDD.n33 95.5247
R166 VDD.n61 VDD.n12 84.8808
R167 VDD.n67 VDD.n66 84.8808
R168 VDD.n62 VDD.t40 81.9927
R169 VDD.n62 VDD.t43 81.9927
R170 VDD.n59 VDD.n57 59.7112
R171 VDD.n68 VDD.n7 57.051
R172 VDD.n37 VDD.n34 55.1976
R173 VDD.n59 VDD.n58 44.8005
R174 VDD.n58 VDD.n7 44.8005
R175 VDD.n41 VDD.n34 34.6747
R176 VDD.n55 VDD.n9 30.8338
R177 VDD.t40 VDD.n9 30.8338
R178 VDD.n65 VDD.n6 30.8338
R179 VDD.n8 VDD.n7 30.8338
R180 VDD.t43 VDD.n8 30.8338
R181 VDD.n60 VDD.n59 30.8338
R182 VDD.n41 VDD.n40 30.8338
R183 VDD.n38 VDD.n37 30.8338
R184 VDD.n61 VDD.n60 30.2553
R185 VDD.n66 VDD.n65 30.2553
R186 VDD.n14 VDD.t13 28.5655
R187 VDD.n14 VDD.t29 28.5655
R188 VDD.n22 VDD.t33 28.5655
R189 VDD.n22 VDD.t37 28.5655
R190 VDD.n21 VDD.t31 28.5655
R191 VDD.n21 VDD.t3 28.5655
R192 VDD.n20 VDD.t19 28.5655
R193 VDD.n20 VDD.t1 28.5655
R194 VDD.n19 VDD.t5 28.5655
R195 VDD.n19 VDD.t25 28.5655
R196 VDD.n18 VDD.t23 28.5655
R197 VDD.n18 VDD.t15 28.5655
R198 VDD.n17 VDD.t21 28.5655
R199 VDD.n17 VDD.t11 28.5655
R200 VDD.n16 VDD.t7 28.5655
R201 VDD.n16 VDD.t39 28.5655
R202 VDD.n15 VDD.t27 28.5655
R203 VDD.n15 VDD.t35 28.5655
R204 VDD.n23 VDD.t9 28.5655
R205 VDD.n23 VDD.t17 28.5655
R206 VDD.n2 VDD.t52 28.5655
R207 VDD.n2 VDD.t44 28.5655
R208 VDD.n0 VDD.t45 28.5655
R209 VDD.n0 VDD.t51 28.5655
R210 VDD.n48 VDD.t48 28.5655
R211 VDD.n48 VDD.t49 28.5655
R212 VDD.n46 VDD.t41 28.5655
R213 VDD.n46 VDD.t47 28.5655
R214 VDD.n42 VDD.n33 16.8245
R215 VDD.n69 VDD.n6 11.9734
R216 VDD.n69 VDD.n68 11.5786
R217 VDD.n56 VDD.n55 10.2507
R218 VDD.n42 VDD.n41 7.47279
R219 VDD.n43 VDD.n42 7.29386
R220 VDD.n55 VDD.n54 6.70286
R221 VDD.n54 VDD.n6 6.70286
R222 VDD.n68 VDD.n67 4.5127
R223 VDD.n63 VDD.n11 4.5127
R224 VDD.n63 VDD.n62 4.5127
R225 VDD.n57 VDD.n12 4.5127
R226 VDD.n35 VDD.n34 3.85467
R227 VDD.n39 VDD.n35 3.85467
R228 VDD.n36 VDD.n33 3.85467
R229 VDD.n39 VDD.n36 3.85467
R230 VDD.n50 VDD.n49 3.44938
R231 VDD.n4 VDD.n3 3.4375
R232 VDD.n43 VDD.n13 2.76114
R233 VDD.n57 VDD.n56 2.72315
R234 VDD.n56 VDD.n53 0.989058
R235 VDD.n53 VDD.n13 0.776701
R236 VDD.n44 VDD.n32 0.525141
R237 VDD.t40 VDD.n61 0.427897
R238 VDD.n66 VDD.t43 0.427897
R239 VDD.n49 VDD.n47 0.239156
R240 VDD.n3 VDD.n1 0.229
R241 VDD.n26 VDD.n25 0.196578
R242 VDD.n28 VDD.n27 0.195966
R243 VDD.n31 VDD.n30 0.195353
R244 VDD.n25 VDD.n24 0.193515
R245 VDD.n30 VDD.n29 0.192902
R246 VDD.n29 VDD.n28 0.192902
R247 VDD.n27 VDD.n26 0.192902
R248 VDD.n52 VDD.n51 0.175096
R249 VDD.n51 VDD.n5 0.160189
R250 VDD.n32 VDD.n31 0.130263
R251 VDD.n70 VDD.n5 0.12602
R252 VDD.n5 VDD.n4 0.061504
R253 VDD.n53 VDD.n52 0.0572073
R254 VDD.n51 VDD.n50 0.0563511
R255 VDD.n45 VDD.n44 0.0502099
R256 VDD.n70 VDD.n69 0.0481923
R257 VDD.n44 VDD.n43 0.0463128
R258 VDD.n45 VDD.n13 0.0397405
R259 VDD VDD.n70 0.0244618
R260 VDD.n52 VDD.n45 0.0144768
R261 VBIAS.t3 VBIAS.n7 50.938
R262 VBIAS.n9 VBIAS.t3 50.938
R263 VBIAS.n6 VBIAS.t5 50.938
R264 VBIAS.t5 VBIAS.n4 50.938
R265 VBIAS.n0 VBIAS.t6 26.3192
R266 VBIAS.n8 VBIAS.t0 25.9322
R267 VBIAS.n5 VBIAS.t7 25.9164
R268 VBIAS.n2 VBIAS.t8 25.6066
R269 VBIAS.n1 VBIAS.t9 25.5864
R270 VBIAS.n0 VBIAS.t10 25.5841
R271 VBIAS.n11 VBIAS.t1 25.3038
R272 VBIAS.n16 VBIAS.t4 25.3038
R273 VBIAS.n13 VBIAS.t2 25.2968
R274 VBIAS.n19 VBIAS.n18 3.12666
R275 VBIAS.n10 VBIAS.n3 1.3304
R276 VBIAS.n15 VBIAS.n6 1.22993
R277 VBIAS.n14 VBIAS.n12 1.21906
R278 VBIAS.n12 VBIAS.n7 1.19188
R279 VBIAS.n17 VBIAS.n4 1.17793
R280 VBIAS.n15 VBIAS.n14 1.17558
R281 VBIAS.n10 VBIAS.n9 1.13989
R282 VBIAS.n18 VBIAS.n17 0.958326
R283 VBIAS.n1 VBIAS.n0 0.717709
R284 VBIAS.n2 VBIAS.n1 0.670292
R285 VBIAS VBIAS.n19 0.566284
R286 VBIAS.n18 VBIAS.n3 0.365632
R287 VBIAS.n13 VBIAS.n3 0.346964
R288 VBIAS.n14 VBIAS.n13 0.346964
R289 VBIAS.n11 VBIAS.n10 0.332875
R290 VBIAS.n12 VBIAS.n11 0.332875
R291 VBIAS.n17 VBIAS.n16 0.332875
R292 VBIAS.n16 VBIAS.n15 0.332875
R293 VBIAS.n8 VBIAS.n7 0.279857
R294 VBIAS.n6 VBIAS.n5 0.278875
R295 VBIAS.n9 VBIAS.n8 0.270541
R296 VBIAS.n5 VBIAS.n4 0.269393
R297 VBIAS.n19 VBIAS.n2 0.148833
R298 VSS.n56 VSS.n5 29835.6
R299 VSS.n57 VSS.n56 23778.9
R300 VSS.n54 VSS.n6 11339.1
R301 VSS.n27 VSS.n6 11339.1
R302 VSS.n54 VSS.n7 11339.1
R303 VSS.n27 VSS.n7 11339.1
R304 VSS.n59 VSS.n2 7358.53
R305 VSS.n59 VSS.n3 6572.62
R306 VSS.n4 VSS.n2 6463.34
R307 VSS.n4 VSS.n3 3664.89
R308 VSS.n56 VSS.n55 3434.98
R309 VSS.n49 VSS.n12 3377.97
R310 VSS.n49 VSS.n13 3377.97
R311 VSS.n40 VSS.n36 3377.97
R312 VSS.n41 VSS.n36 3377.97
R313 VSS.n48 VSS.n29 2297.58
R314 VSS.n45 VSS.n30 2259.71
R315 VSS.n45 VSS.n31 2259.71
R316 VSS.n30 VSS.n12 1118.26
R317 VSS.n40 VSS.n30 1118.26
R318 VSS.n31 VSS.n13 1118.26
R319 VSS.n41 VSS.n31 1118.26
R320 VSS.t13 VSS.t18 922.712
R321 VSS.t16 VSS.t13 922.712
R322 VSS.n53 VSS.n8 736.754
R323 VSS.n53 VSS.n52 732.236
R324 VSS.t7 VSS.n3 725.548
R325 VSS.n55 VSS.t18 691.027
R326 VSS.n29 VSS.t16 676.923
R327 VSS.t3 VSS.n5 455.969
R328 VSS.t5 VSS.n57 447.098
R329 VSS.n58 VSS.t1 406.291
R330 VSS.n58 VSS.t5 406.291
R331 VSS.n57 VSS.t7 365.485
R332 VSS.t20 VSS.n46 342.42
R333 VSS.t0 VSS.n37 342.42
R334 VSS.t0 VSS.t10 312.259
R335 VSS.n47 VSS.t20 235.969
R336 VSS.n42 VSS.n41 195
R337 VSS.n41 VSS.t0 195
R338 VSS.n35 VSS.n13 195
R339 VSS.t20 VSS.n13 195
R340 VSS.n12 VSS.n11 195
R341 VSS.t20 VSS.n12 195
R342 VSS.n40 VSS.n39 195
R343 VSS.t0 VSS.n40 195
R344 VSS.n25 VSS.n8 187.482
R345 VSS.n37 VSS.t1 157.904
R346 VSS.n44 VSS.n32 146.825
R347 VSS.n44 VSS.n43 146.825
R348 VSS.n28 VSS.t3 123.246
R349 VSS.n3 VSS.n1 117.001
R350 VSS.n27 VSS.n26 117.001
R351 VSS.t3 VSS.n27 117.001
R352 VSS.n10 VSS.n2 117.001
R353 VSS.n47 VSS.n2 117.001
R354 VSS.n54 VSS.n53 117.001
R355 VSS.n55 VSS.n54 117.001
R356 VSS.n28 VSS.n7 116.275
R357 VSS.n48 VSS.n47 106.453
R358 VSS.n21 VSS.t8 86.18
R359 VSS.n20 VSS.t11 86.1487
R360 VSS.n24 VSS.t9 83.7172
R361 VSS.n32 VSS.n11 72.6593
R362 VSS.n39 VSS.n32 72.6593
R363 VSS.n33 VSS.n1 71.3578
R364 VSS.n39 VSS.n38 69.9281
R365 VSS.n16 VSS.n14 69.7168
R366 VSS.n18 VSS.n17 69.5228
R367 VSS.n16 VSS.n15 69.5222
R368 VSS.n20 VSS.n19 68.2652
R369 VSS.n50 VSS.n11 66.5266
R370 VSS.n45 VSS.n44 58.5005
R371 VSS.n46 VSS.n45 58.5005
R372 VSS.n38 VSS.n36 58.5005
R373 VSS.n37 VSS.n36 58.5005
R374 VSS.n50 VSS.n49 58.5005
R375 VSS.n49 VSS.n48 58.5005
R376 VSS.n29 VSS.n28 56.1087
R377 VSS.n60 VSS.n1 42.8204
R378 VSS.n46 VSS.t10 30.1618
R379 VSS.n34 VSS.n33 27.7065
R380 VSS.n33 VSS.n4 20.8934
R381 VSS.n58 VSS.n4 20.8934
R382 VSS.n60 VSS.n59 20.8934
R383 VSS.n59 VSS.n58 20.8934
R384 VSS.n19 VSS.t2 17.4005
R385 VSS.n19 VSS.t6 17.4005
R386 VSS.n14 VSS.t19 17.4005
R387 VSS.n14 VSS.t14 17.4005
R388 VSS.n15 VSS.t17 17.4005
R389 VSS.n15 VSS.t15 17.4005
R390 VSS.n17 VSS.t12 17.4005
R391 VSS.n17 VSS.t4 17.4005
R392 VSS.n52 VSS.n7 12.188
R393 VSS.n8 VSS.n6 12.188
R394 VSS.n6 VSS.n5 12.188
R395 VSS.n52 VSS.n51 11.1022
R396 VSS.n51 VSS.n50 11.1022
R397 VSS.n26 VSS.n9 8.97973
R398 VSS.n51 VSS.n10 6.30179
R399 VSS.n38 VSS.n0 6.25627
R400 VSS.n26 VSS.n25 4.78618
R401 VSS.n43 VSS.n35 4.06366
R402 VSS.n43 VSS.n42 4.06366
R403 VSS.n42 VSS.n0 3.70576
R404 VSS.n24 VSS.n18 3.39902
R405 VSS.n25 VSS.n24 3.15791
R406 VSS.n35 VSS.n34 2.44261
R407 VSS.n51 VSS.n9 1.63752
R408 VSS VSS.n0 1.62304
R409 VSS VSS.n60 0.965007
R410 VSS.n23 VSS.n22 0.504422
R411 VSS.n22 VSS 0.328244
R412 VSS.n18 VSS.n16 0.192906
R413 VSS.n24 VSS.n23 0.148333
R414 VSS.n34 VSS.n10 0.140346
R415 VSS.n22 VSS.n21 0.0780862
R416 VSS.n23 VSS.n9 0.0299304
R417 VSS.n21 VSS.n20 0.00101653
R418 V2.n0 V2.n4 199.65
R419 V2.t3 V2.n0 25.9937
R420 V2.n0 V2.t11 25.8614
R421 V2.t9 V2.n1 25.8883
R422 V2.n0 V2.t5 25.8406
R423 V2.t7 V2.n0 25.9857
R424 V2.n0 V2.t0 35.7682
R425 V2.n4 V2.t6 28.5655
R426 V2.n4 V2.t8 28.5655
R427 V2.n3 V2.t12 28.5655
R428 V2.n3 V2.t10 28.5655
R429 V2.n2 V2.t2 28.5655
R430 V2.n2 V2.t4 28.5655
R431 V2.n0 V2.t13 26.2697
R432 V2.n0 V2.t16 26.2675
R433 V2.n0 V2.t18 26.2568
R434 V2.n0 V2.t14 26.2558
R435 V2.n0 V2.t17 26.2556
R436 V2.n0 V2.t15 26.2553
R437 V2.n1 V2.n0 0.249974
R438 V2.n0 V2.t1 26.0106
R439 V2.n0 V2.n2 200.287
R440 V2.n1 V2.n3 199.899
R441 MINUS MINUS.t0 161.175
R442 PLUS PLUS.t0 157.964
C0 VDD MINUS 0.015211f
C1 PLUS MINUS 0.356659f
C2 VOUT V1 2.01272f
C3 a_2586_n2492# MINUS 0.566541f
C4 PLUS VDD 0.032248f
C5 VBIAS VOUT 2.09473f
C6 a_2586_n2492# VDD 0.068018f
C7 PLUS a_2586_n2492# 0.345141f
C8 VOUT VDD 7.55246f
C9 VBIAS V1 0.198595f
C10 PLUS VOUT 0.022003f
C11 V1 MINUS 0.02059f
C12 VBIAS MINUS 0.603904f
C13 V1 VDD 11.3658f
C14 PLUS V1 0.388481f
C15 V1 a_2586_n2492# 0.108067f
C16 VBIAS VDD 0.338353f
C17 VBIAS PLUS 0.458357f
C18 VBIAS a_2586_n2492# 1.43327f
.ends

