magic
tech sky130A
timestamp 1713067979
<< pwell >>
rect -341 -489 341 489
<< nmos >>
rect -243 -384 -143 415
rect -114 -384 -14 415
rect 14 -384 114 415
rect 143 -384 243 415
<< ndiff >>
rect -272 409 -243 415
rect -272 -378 -266 409
rect -249 -378 -243 409
rect -272 -384 -243 -378
rect -143 409 -114 415
rect -143 -378 -137 409
rect -120 -378 -114 409
rect -143 -384 -114 -378
rect -14 409 14 415
rect -14 -378 -8 409
rect 8 -378 14 409
rect -14 -384 14 -378
rect 114 409 143 415
rect 114 -378 120 409
rect 137 -378 143 409
rect 114 -384 143 -378
rect 243 409 272 415
rect 243 -378 249 409
rect 266 -378 272 409
rect 243 -384 272 -378
<< ndiffc >>
rect -266 -378 -249 409
rect -137 -378 -120 409
rect -8 -378 8 409
rect 120 -378 137 409
rect 249 -378 266 409
<< psubdiff >>
rect -323 454 323 471
rect -323 423 -306 454
rect 306 423 323 454
rect -323 -454 -306 -423
rect 306 -454 323 -423
rect -323 -471 -275 -454
rect 275 -471 323 -454
<< psubdiffcont >>
rect -323 -423 -306 423
rect 306 -423 323 423
rect -275 -471 275 -454
<< poly >>
rect -243 415 -143 428
rect -114 415 -14 428
rect 14 415 114 428
rect 143 415 243 428
rect -243 -403 -143 -384
rect -243 -420 -235 -403
rect -151 -420 -143 -403
rect -243 -428 -143 -420
rect -114 -403 -14 -384
rect -114 -420 -106 -403
rect -22 -420 -14 -403
rect -114 -428 -14 -420
rect 14 -403 114 -384
rect 14 -420 22 -403
rect 106 -420 114 -403
rect 14 -428 114 -420
rect 143 -403 243 -384
rect 143 -420 151 -403
rect 235 -420 243 -403
rect 143 -428 243 -420
<< polycont >>
rect -235 -420 -151 -403
rect -106 -420 -22 -403
rect 22 -420 106 -403
rect 151 -420 235 -403
<< locali >>
rect -323 423 -306 471
rect 306 423 323 471
rect -266 409 -249 417
rect -266 -386 -249 -378
rect -137 409 -120 417
rect -137 -386 -120 -378
rect -8 409 8 417
rect -8 -386 8 -378
rect 120 409 137 417
rect 120 -386 137 -378
rect 249 409 266 417
rect 249 -386 266 -378
rect -243 -420 -235 -403
rect -151 -420 -143 -403
rect -114 -420 -106 -403
rect -22 -420 -14 -403
rect 14 -420 22 -403
rect 106 -420 114 -403
rect 143 -420 151 -403
rect 235 -420 243 -403
rect -323 -471 -275 -454
rect 275 -471 323 -454
<< viali >>
rect -306 454 306 471
rect -323 -423 -306 -91
rect -266 86 -249 401
rect -137 -370 -120 -55
rect -8 86 8 401
rect 120 -370 137 -55
rect 249 86 266 401
rect -235 -420 -151 -403
rect -106 -420 -22 -403
rect 22 -420 106 -403
rect 151 -420 235 -403
rect -323 -454 -306 -423
rect 306 -423 323 -91
rect 306 -454 323 -423
<< metal1 >>
rect -312 471 312 474
rect -312 454 -306 471
rect 306 454 312 471
rect -312 451 312 454
rect -269 401 -246 407
rect -269 86 -266 401
rect -249 86 -246 401
rect -269 80 -246 86
rect -11 401 11 407
rect -11 86 -8 401
rect 8 86 11 401
rect -11 80 11 86
rect 246 401 269 407
rect 246 86 249 401
rect 266 86 269 401
rect 246 80 269 86
rect -140 -55 -117 -49
rect -326 -91 -303 -85
rect -326 -454 -323 -91
rect -306 -454 -303 -91
rect -140 -370 -137 -55
rect -120 -370 -117 -55
rect -140 -376 -117 -370
rect 117 -55 140 -49
rect 117 -370 120 -55
rect 137 -370 140 -55
rect 117 -376 140 -370
rect 303 -91 326 -85
rect -241 -403 -145 -400
rect -241 -420 -235 -403
rect -151 -420 -145 -403
rect -241 -423 -145 -420
rect -112 -403 -16 -400
rect -112 -420 -106 -403
rect -22 -420 -16 -403
rect -112 -423 -16 -420
rect 16 -403 112 -400
rect 16 -420 22 -403
rect 106 -420 112 -403
rect 16 -423 112 -420
rect 145 -403 241 -400
rect 145 -420 151 -403
rect 235 -420 241 -403
rect 145 -423 241 -420
rect -326 -460 -303 -454
rect 303 -454 306 -91
rect 323 -454 326 -91
rect 303 -460 326 -454
<< properties >>
string FIXED_BBOX -315 -463 315 463
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
