magic
tech sky130A
magscale 1 2
timestamp 1713539272
<< pwell >>
rect -425 -3410 425 3410
<< nmoslvt >>
rect -229 -3200 -29 3200
rect 29 -3200 229 3200
<< ndiff >>
rect -287 3188 -229 3200
rect -287 -3188 -275 3188
rect -241 -3188 -229 3188
rect -287 -3200 -229 -3188
rect -29 3188 29 3200
rect -29 -3188 -17 3188
rect 17 -3188 29 3188
rect -29 -3200 29 -3188
rect 229 3188 287 3200
rect 229 -3188 241 3188
rect 275 -3188 287 3188
rect 229 -3200 287 -3188
<< ndiffc >>
rect -275 -3188 -241 3188
rect -17 -3188 17 3188
rect 241 -3188 275 3188
<< psubdiff >>
rect -389 3340 -293 3374
rect 293 3340 389 3374
rect -389 3278 -355 3340
rect 355 3278 389 3340
rect -389 -3340 -355 -3278
rect 355 -3340 389 -3278
rect -389 -3374 -293 -3340
rect 293 -3374 389 -3340
<< psubdiffcont >>
rect -293 3340 293 3374
rect -389 -3278 -355 3278
rect 355 -3278 389 3278
rect -293 -3374 293 -3340
<< poly >>
rect -229 3272 -29 3288
rect -229 3238 -213 3272
rect -45 3238 -29 3272
rect -229 3200 -29 3238
rect 29 3272 229 3288
rect 29 3238 45 3272
rect 213 3238 229 3272
rect 29 3200 229 3238
rect -229 -3238 -29 -3200
rect -229 -3272 -213 -3238
rect -45 -3272 -29 -3238
rect -229 -3288 -29 -3272
rect 29 -3238 229 -3200
rect 29 -3272 45 -3238
rect 213 -3272 229 -3238
rect 29 -3288 229 -3272
<< polycont >>
rect -213 3238 -45 3272
rect 45 3238 213 3272
rect -213 -3272 -45 -3238
rect 45 -3272 213 -3238
<< locali >>
rect -389 3340 -293 3374
rect 293 3340 389 3374
rect -389 3278 -355 3340
rect 355 3278 389 3340
rect -229 3238 -213 3272
rect -45 3238 -29 3272
rect 29 3238 45 3272
rect 213 3238 229 3272
rect -275 3188 -241 3204
rect -275 -3204 -241 -3188
rect -17 3188 17 3204
rect -17 -3204 17 -3188
rect 241 3188 275 3204
rect 241 -3204 275 -3188
rect -229 -3272 -213 -3238
rect -45 -3272 -29 -3238
rect 29 -3272 45 -3238
rect 213 -3272 229 -3238
rect -389 -3340 -355 -3278
rect 355 -3340 389 -3278
rect -389 -3374 -293 -3340
rect 293 -3374 389 -3340
<< viali >>
rect -213 3238 -45 3272
rect 45 3238 213 3272
rect -275 -3188 -241 3188
rect -17 -3188 17 3188
rect 241 -3188 275 3188
rect -213 -3272 -45 -3238
rect 45 -3272 213 -3238
<< metal1 >>
rect -225 3272 -33 3278
rect -225 3238 -213 3272
rect -45 3238 -33 3272
rect -225 3232 -33 3238
rect 33 3272 225 3278
rect 33 3238 45 3272
rect 213 3238 225 3272
rect 33 3232 225 3238
rect -281 3188 -235 3200
rect -281 -3188 -275 3188
rect -241 -3188 -235 3188
rect -281 -3200 -235 -3188
rect -23 3188 23 3200
rect -23 -3188 -17 3188
rect 17 -3188 23 3188
rect -23 -3200 23 -3188
rect 235 3188 281 3200
rect 235 -3188 241 3188
rect 275 -3188 281 3188
rect 235 -3200 281 -3188
rect -225 -3238 -33 -3232
rect -225 -3272 -213 -3238
rect -45 -3272 -33 -3238
rect -225 -3278 -33 -3272
rect 33 -3238 225 -3232
rect 33 -3272 45 -3238
rect 213 -3272 225 -3238
rect 33 -3278 225 -3272
<< properties >>
string FIXED_BBOX -372 -3357 372 3357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 32.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
