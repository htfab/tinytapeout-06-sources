magic
tech sky130A
magscale 1 2
timestamp 1713550165
<< pwell >>
rect 40 2200 140 2600
rect 560 2580 620 2740
rect 1460 -330 1480 3080
rect 1500 3040 1570 3130
rect 3000 -120 3080 560
rect 4510 -120 4520 530
rect 3000 -160 3580 -120
rect 4070 -140 4130 -120
rect 3000 -200 3040 -160
rect 3132 -164 3460 -160
<< nmoslvt >>
rect 40 2200 140 2600
rect 560 2580 620 2740
<< locali >>
rect -1000 10200 6600 10400
rect -1000 9880 -690 10200
rect 6300 9880 6600 10200
rect -1000 9800 6600 9880
rect -1000 9700 5400 9800
rect -1000 7700 -500 9700
rect -100 7700 300 9700
rect 700 7700 900 9700
rect 1300 9640 5400 9700
rect 1300 9600 5390 9640
rect 1300 7700 1600 9600
rect -1000 7400 1600 7700
rect -1000 6000 -400 7400
rect 400 6000 600 7400
rect 1200 6000 1600 7400
rect 2600 6000 2800 9600
rect 3800 6000 4000 9600
rect 5000 6300 5100 9600
rect 5300 6300 5390 9600
rect 5000 6000 5390 6300
rect -1000 5584 3260 5640
rect -1000 5550 -268 5584
rect 60 5550 532 5584
rect 860 5550 3260 5584
rect -1000 5540 3260 5550
rect -1000 5500 -280 5540
rect 80 5500 440 5540
rect -1000 5488 -340 5500
rect 130 5488 440 5500
rect 920 5536 1460 5540
rect -1000 3732 -364 5488
rect 130 3732 436 5488
rect 954 5488 1460 5536
rect 1940 5488 2260 5540
rect 954 3780 1436 5488
rect 920 3732 1436 3780
rect 1956 3732 2236 5488
rect -1000 3660 -340 3732
rect 130 3660 440 3732
rect 920 3660 1460 3732
rect 1940 3660 2260 3732
rect 2720 3660 3200 5540
rect -1000 3180 3200 3660
rect -1000 3126 -360 3180
rect -1000 -230 -400 3126
rect -366 -230 -360 3126
rect 840 3130 3200 3180
rect 840 3126 1500 3130
rect -1000 -290 -360 -230
rect 840 -230 860 3126
rect 894 3088 1500 3126
rect 894 -230 1436 3088
rect 840 -268 1436 -230
rect 1470 -268 1500 3088
rect 2700 2000 3200 3130
rect 3800 2000 4000 5600
rect 4800 2210 5390 5600
rect 4800 2190 5710 2210
rect 4800 2000 6600 2190
rect 2700 1720 6600 2000
rect 2700 1480 3070 1720
rect 6080 1480 6600 1720
rect 2700 1130 6600 1480
rect 2700 870 3070 1130
rect 6080 870 6600 1130
rect 2700 584 6600 870
rect 2700 550 3132 584
rect 3460 550 4132 584
rect 4460 550 6600 584
rect 2700 -30 3080 550
rect 3500 540 6600 550
rect 3500 488 4080 540
rect 3500 390 3522 488
rect 3442 22 3522 390
rect 2700 -68 3036 -30
rect 3070 -68 3080 -30
rect 2700 -120 3080 -68
rect 3500 -68 3522 22
rect 3556 -68 4036 488
rect 4070 -68 4080 488
rect 4210 482 4380 500
rect 4460 490 6600 540
rect 4540 488 6600 490
rect 4210 448 4212 482
rect 4210 440 4380 448
rect 4230 430 4370 440
rect 4300 290 4370 430
rect 4184 90 4370 290
rect 4300 -10 4370 90
rect 4442 40 4522 380
rect 4230 -20 4370 -10
rect 3500 -120 4080 -68
rect 4210 -28 4380 -20
rect 4210 -62 4212 -28
rect 4210 -80 4380 -62
rect 4490 -68 4522 -60
rect 4556 -68 6600 488
rect 4490 -90 6600 -68
rect 2700 -130 4130 -120
rect 2700 -164 3132 -130
rect 3460 -164 4132 -130
rect 4460 -164 6600 -90
rect 840 -290 1500 -268
rect -1000 -330 1500 -290
rect 2700 -330 6600 -164
rect -1000 -1000 6600 -330
<< viali >>
rect -690 9880 6300 10200
rect -500 7700 -100 9700
rect 300 7700 700 9700
rect 900 7700 1300 9700
rect 5100 6300 5300 9600
rect -268 5550 60 5584
rect 532 5550 860 5584
rect -364 3732 -330 5488
rect -188 5448 -20 5482
rect -250 3822 -216 5398
rect 436 3732 470 5488
rect 920 3780 954 5536
rect 1436 3732 1470 5488
rect 1922 3732 1956 5488
rect 2236 3732 2270 5488
rect -400 -230 -366 3126
rect -286 -140 -252 3036
rect -28 -140 6 3036
rect 230 -140 264 3036
rect 488 -140 522 3036
rect 746 -140 780 3036
rect -224 -224 -56 -190
rect 34 -224 202 -190
rect 292 -224 460 -190
rect 550 -224 718 -190
rect 860 -230 894 3126
rect 1436 -268 1470 3088
rect 5566 1566 5998 1636
rect 3166 966 3598 1036
rect 5566 966 5998 1036
rect 3132 550 3460 584
rect 4132 550 4460 584
rect 3212 448 3380 482
rect 3150 22 3184 398
rect 3408 22 3442 398
rect 3036 -68 3070 -30
rect 3212 -62 3380 -28
rect 3522 -68 3556 488
rect 4036 -68 4070 488
rect 4212 448 4380 482
rect 4150 22 4184 398
rect 4408 22 4442 398
rect 4212 -62 4380 -28
rect 4522 -68 4556 488
rect 3132 -164 3460 -130
rect 4132 -164 4460 -130
rect 1612 -262 1780 -228
rect 1870 -262 2038 -228
rect 2128 -262 2296 -228
rect 2386 -262 2554 -228
<< metal1 >>
rect -1000 10200 6600 10400
rect -1000 9880 -690 10200
rect 6300 9880 6600 10200
rect -1000 9800 6600 9880
rect -1000 9700 5400 9800
rect -1000 7700 -500 9700
rect -100 7700 300 9700
rect 700 7700 900 9700
rect 1300 9640 5400 9700
rect 1300 9600 5390 9640
rect 1300 7700 1600 9600
rect -1000 7400 1600 7700
rect -1000 6000 -400 7400
rect 400 6000 600 7400
rect 1200 6000 1600 7400
rect 2600 6000 2800 9600
rect 3800 6000 4000 9600
rect 5000 6300 5100 9600
rect 5300 6300 5390 9600
rect 5000 6000 5390 6300
rect -1000 5584 3260 5640
rect -1000 5550 -268 5584
rect 60 5550 532 5584
rect 860 5550 3260 5584
rect -1000 5540 3260 5550
rect -1000 5500 -280 5540
rect 80 5500 440 5540
rect 914 5536 1460 5540
rect -1000 5488 -324 5500
rect 130 5488 476 5500
rect -1000 3732 -364 5488
rect -330 3732 -324 5488
rect -200 5482 -8 5488
rect -200 5448 -188 5482
rect -20 5448 -8 5482
rect -200 5442 -8 5448
rect -256 5398 -210 5410
rect -256 3822 -250 5398
rect -216 5040 -210 5398
rect -180 5140 -40 5442
rect -160 4920 -150 5040
rect -216 3822 -210 4920
rect -120 4880 -40 5140
rect -256 3810 -210 3822
rect -180 4760 -40 4880
rect -180 4640 -150 4760
rect -70 4640 -40 4760
rect -180 3740 -40 4640
rect -10 4040 0 4120
rect 80 4040 90 4120
rect -1000 3720 -324 3732
rect 130 3732 436 5488
rect 470 3732 476 5488
rect 630 5400 770 5480
rect 630 5200 740 5400
rect 790 5220 800 5380
rect 860 5220 870 5380
rect 630 4450 770 5200
rect 630 4330 660 4450
rect 740 4330 770 4450
rect 630 4180 770 4330
rect 530 4040 540 4120
rect 620 4040 630 4120
rect 660 3980 770 4180
rect 630 3740 770 3980
rect 914 3780 920 5536
rect 954 5500 1460 5536
rect 1940 5500 2260 5540
rect 954 5488 1476 5500
rect 954 3780 1436 5488
rect 914 3768 1436 3780
rect 130 3720 476 3732
rect 920 3732 1436 3768
rect 1470 3732 1476 5488
rect 1916 5488 2276 5500
rect 1630 5140 1770 5480
rect 1530 4900 1540 5100
rect 1600 4900 1610 5100
rect 1660 4860 1770 5140
rect 1630 4460 1770 4860
rect 1630 4340 1660 4460
rect 1740 4340 1770 4460
rect 1630 4200 1770 4340
rect 1630 3960 1720 4200
rect 1760 4020 1780 4100
rect 1840 4020 1850 4100
rect 1630 3740 1770 3960
rect 920 3720 1476 3732
rect 1916 3732 1922 5488
rect 1956 3732 2236 5488
rect 2270 3732 2276 5488
rect 2430 5400 2570 5490
rect 2430 5180 2560 5400
rect 2590 5200 2600 5380
rect 2660 5200 2670 5380
rect 2430 4750 2570 5180
rect 2430 4630 2450 4750
rect 2530 4630 2570 4750
rect 2430 4240 2570 4630
rect 2350 4020 2360 4100
rect 2440 4020 2450 4100
rect 2480 3940 2570 4240
rect 2430 3750 2570 3940
rect 1916 3720 2276 3732
rect -1000 3660 -340 3720
rect 130 3660 440 3720
rect 920 3660 1460 3720
rect 1940 3660 2260 3720
rect 2720 3660 3200 5540
rect -1000 3180 3200 3660
rect -1000 3126 -360 3180
rect -1000 -230 -400 3126
rect -366 -230 -360 3126
rect 850 3130 3200 3180
rect 850 3126 1500 3130
rect -292 3036 -246 3048
rect -292 2540 -286 3036
rect -300 2300 -286 2540
rect -252 2540 -246 3036
rect -190 2560 -106 3114
rect -252 2480 -210 2540
rect -292 -140 -286 2300
rect -252 2300 -210 2320
rect -252 -140 -246 2300
rect -170 2250 -106 2560
rect -292 -152 -246 -140
rect -190 1500 -106 2250
rect -190 1380 -180 1500
rect -120 1380 -106 1500
rect -190 -184 -106 1380
rect -34 3036 12 3048
rect -34 250 -28 3036
rect 6 250 12 3036
rect 80 2620 164 3104
rect 224 3036 270 3048
rect 80 2600 140 2620
rect 40 2220 140 2600
rect 224 2480 230 3036
rect 264 2480 270 3036
rect 320 2560 404 3114
rect 482 3036 528 3048
rect 320 2520 420 2560
rect 190 2340 200 2480
rect 300 2340 310 2480
rect 40 2200 164 2220
rect 80 1500 164 2200
rect 80 1380 100 1500
rect 160 1380 170 1500
rect -70 100 -60 250
rect 40 100 50 250
rect -34 -140 -28 100
rect 6 -140 12 100
rect -34 -152 12 -140
rect 80 -184 164 1380
rect 224 -140 230 2340
rect 264 -140 270 2340
rect 340 2300 420 2520
rect 224 -152 270 -140
rect 320 2280 420 2300
rect 320 1520 404 2280
rect 320 1400 340 1520
rect 400 1400 410 1520
rect 320 290 404 1400
rect 320 90 390 290
rect 482 250 488 3036
rect 522 250 528 3036
rect 600 2880 684 3094
rect 560 2760 684 2880
rect 740 3036 786 3048
rect 560 2480 640 2760
rect 740 2540 746 3036
rect 780 2540 786 3036
rect 560 2300 620 2480
rect 690 2340 700 2540
rect 780 2340 790 2540
rect 560 2220 640 2300
rect 560 2180 684 2220
rect 580 2040 684 2180
rect 600 1500 684 2040
rect 600 1380 620 1500
rect 680 1380 690 1500
rect 430 120 450 250
rect 560 120 570 250
rect 320 -184 404 90
rect 482 -140 488 120
rect 522 -140 528 120
rect 482 -152 528 -140
rect 600 -184 684 1380
rect 740 -140 746 2340
rect 780 -140 786 2340
rect 740 -152 786 -140
rect -236 -190 -44 -184
rect -236 -224 -224 -190
rect -56 -224 -44 -190
rect -236 -230 -44 -224
rect 22 -190 214 -184
rect 22 -224 34 -190
rect 202 -224 214 -190
rect 22 -230 214 -224
rect 280 -190 472 -184
rect 280 -224 292 -190
rect 460 -224 472 -190
rect 280 -230 472 -224
rect 538 -190 730 -184
rect 538 -224 550 -190
rect 718 -224 730 -190
rect 538 -230 730 -224
rect 850 -230 860 3126
rect 894 3088 1500 3126
rect 894 -230 1436 3088
rect -1000 -290 -360 -230
rect 850 -268 1436 -230
rect 1470 3050 1500 3088
rect 1470 -268 1480 3050
rect 1640 2650 1724 3074
rect 1640 2640 1760 2650
rect 1650 2360 1660 2560
rect 1690 2290 1760 2640
rect 1690 2280 1724 2290
rect 1640 900 1724 2280
rect 1920 920 2000 3070
rect 2030 2340 2040 2540
rect 2120 2340 2130 2540
rect 2170 920 2250 3090
rect 1640 780 1660 900
rect 1720 780 1730 900
rect 1920 800 1940 920
rect 2000 800 2010 920
rect 2170 800 2180 920
rect 2240 800 2250 920
rect 1640 -222 1724 780
rect 1920 300 2000 800
rect 1760 110 1770 240
rect 1890 110 1900 240
rect 1940 50 2000 300
rect 1920 -222 2000 50
rect 2170 -222 2250 800
rect 2440 940 2520 3090
rect 2550 2320 2560 2520
rect 2640 2320 2650 2520
rect 2700 2000 3200 3130
rect 3800 2000 4000 5600
rect 4800 2210 5390 5600
rect 5530 2910 6051 9800
rect 5524 2390 5530 2910
rect 6050 2390 6056 2910
rect 4800 2190 5710 2210
rect 4800 2000 6600 2190
rect 2700 1720 6600 2000
rect 2700 1480 3070 1720
rect 5554 1636 6010 1642
rect 5554 1566 5566 1636
rect 5998 1566 6010 1636
rect 5554 1560 6010 1566
rect 6080 1480 6600 1720
rect 2700 1130 6600 1480
rect 2440 820 2460 940
rect 2520 820 2530 940
rect 2700 870 3070 1130
rect 3154 1036 3610 1042
rect 3154 966 3166 1036
rect 3598 966 3610 1036
rect 3154 960 3610 966
rect 5554 1036 6010 1042
rect 5554 966 5566 1036
rect 5998 966 6010 1036
rect 5554 960 6010 966
rect 6080 870 6600 1130
rect 2440 310 2520 820
rect 2280 130 2290 260
rect 2410 130 2420 260
rect 2460 60 2520 310
rect 2440 -222 2520 60
rect 2700 584 6600 870
rect 2700 550 3132 584
rect 3460 550 4132 584
rect 4460 550 6600 584
rect 2700 -30 3080 550
rect 3120 544 3472 550
rect 3500 540 6600 550
rect 3500 488 4080 540
rect 3200 482 3392 488
rect 3200 448 3212 482
rect 3380 448 3392 482
rect 3200 442 3392 448
rect 3144 400 3190 410
rect 3110 30 3120 400
rect 3180 398 3190 400
rect 3144 22 3150 30
rect 3184 22 3190 398
rect 3144 10 3190 22
rect 3250 300 3340 442
rect 3250 90 3260 300
rect 3320 90 3340 300
rect 3250 -22 3340 90
rect 3402 398 3448 410
rect 3402 22 3408 398
rect 3442 390 3448 398
rect 3500 390 3522 488
rect 3442 22 3522 390
rect 3402 10 3448 22
rect 2700 -68 3036 -30
rect 3070 -68 3080 -30
rect 3200 -28 3392 -22
rect 3200 -62 3212 -28
rect 3380 -62 3392 -28
rect 3200 -68 3392 -62
rect 3500 -68 3522 22
rect 3556 -68 4036 488
rect 4070 -68 4080 488
rect 4150 488 4380 500
rect 4460 490 6600 540
rect 4516 488 6600 490
rect 4150 482 4392 488
rect 4150 448 4212 482
rect 4380 448 4392 482
rect 4150 442 4392 448
rect 4150 440 4380 442
rect 4150 410 4370 440
rect 4144 398 4370 410
rect 4144 22 4150 398
rect 4184 270 4370 398
rect 4402 398 4448 410
rect 4402 380 4408 398
rect 4184 130 4280 270
rect 4340 130 4370 270
rect 4184 22 4370 130
rect 4400 50 4408 380
rect 4144 10 4190 22
rect 4260 -10 4370 22
rect 4402 22 4408 50
rect 4442 380 4448 398
rect 4516 380 4522 488
rect 4442 40 4522 380
rect 4442 22 4448 40
rect 4402 10 4448 22
rect 4230 -20 4370 -10
rect 4210 -22 4380 -20
rect 4200 -28 4380 -22
rect 4200 -62 4212 -28
rect 4516 -60 4522 40
rect 4200 -68 4380 -62
rect 4490 -68 4522 -60
rect 4556 -68 6600 488
rect 2700 -120 3080 -68
rect 3500 -120 4080 -68
rect 4490 -90 6600 -68
rect 2700 -124 3160 -120
rect 3430 -124 4130 -120
rect 4460 -124 6600 -90
rect 2700 -130 6600 -124
rect 2700 -164 3132 -130
rect 3460 -164 4132 -130
rect 4460 -164 6600 -130
rect 1600 -228 1792 -222
rect 1600 -262 1612 -228
rect 1780 -262 1792 -228
rect 1600 -268 1792 -262
rect 1858 -228 2050 -222
rect 1858 -262 1870 -228
rect 2038 -262 2050 -228
rect 1858 -268 2050 -262
rect 2116 -228 2308 -222
rect 2116 -262 2128 -228
rect 2296 -262 2308 -228
rect 2116 -268 2308 -262
rect 2374 -228 2566 -222
rect 2374 -262 2386 -228
rect 2554 -262 2566 -228
rect 2374 -268 2566 -262
rect 850 -290 1480 -268
rect 1920 -270 2000 -268
rect -1000 -330 1480 -290
rect 2700 -330 6600 -164
rect -1000 -1000 6600 -330
<< via1 >>
rect -240 4920 -216 5040
rect -216 4920 -160 5040
rect -150 4640 -70 4760
rect 0 4040 80 4120
rect 800 5220 860 5380
rect 660 4330 740 4450
rect 540 4040 620 4120
rect 1540 4900 1600 5100
rect 1660 4340 1740 4460
rect 1780 4020 1840 4100
rect 2600 5200 2660 5380
rect 2450 4630 2530 4750
rect 2360 4020 2440 4100
rect -280 2320 -252 2480
rect -252 2320 -210 2480
rect -180 1380 -120 1500
rect 200 2340 230 2480
rect 230 2340 264 2480
rect 264 2340 300 2480
rect 100 1380 160 1500
rect -60 100 -28 250
rect -28 100 6 250
rect 6 100 40 250
rect 340 1400 400 1520
rect 700 2340 746 2540
rect 746 2340 780 2540
rect 620 1380 680 1500
rect 450 120 488 250
rect 488 120 522 250
rect 522 120 560 250
rect 1550 2360 1650 2560
rect 2040 2340 2120 2540
rect 1660 780 1720 900
rect 1940 800 2000 920
rect 2180 800 2240 920
rect 1770 110 1890 240
rect 2560 2320 2640 2520
rect 5530 2390 6050 2910
rect 5566 1566 5998 1636
rect 2460 820 2520 940
rect 3166 966 3598 1036
rect 5566 966 5998 1036
rect 2290 130 2410 260
rect 3120 398 3180 400
rect 3120 30 3150 398
rect 3150 30 3180 398
rect 3260 90 3320 300
rect 4280 130 4340 270
<< metal2 >>
rect -1000 5380 3100 5400
rect -1000 5220 800 5380
rect 860 5220 2600 5380
rect -1000 5200 2600 5220
rect 2660 5200 3100 5380
rect 2600 5190 2660 5200
rect 1540 5100 1600 5110
rect -1000 5040 1540 5100
rect -1000 4920 -240 5040
rect -160 4920 1540 5040
rect -1000 4900 1540 4920
rect 1600 4900 3100 5100
rect 1540 4890 1600 4900
rect -1000 4760 3100 4800
rect -1000 4640 -150 4760
rect -70 4750 3100 4760
rect -70 4640 2450 4750
rect -1000 4630 2450 4640
rect 2530 4630 3100 4750
rect -1000 4600 3100 4630
rect -1000 4460 3100 4500
rect -1000 4450 1660 4460
rect -1000 4330 660 4450
rect 740 4340 1660 4450
rect 1740 4340 3100 4460
rect 740 4330 3100 4340
rect -1000 4300 3100 4330
rect -600 4120 1100 4200
rect -600 4040 0 4120
rect 80 4040 540 4120
rect 620 4040 1100 4120
rect -600 4000 1100 4040
rect 1300 4100 3100 4200
rect 1300 4020 1780 4100
rect 1840 4020 2360 4100
rect 2440 4020 3100 4100
rect 1300 4000 3100 4020
rect 100 2700 400 4000
rect 1900 2700 2200 4000
rect 5530 2910 6050 2916
rect -500 2540 1100 2700
rect -500 2480 700 2540
rect -500 2320 -280 2480
rect -210 2340 200 2480
rect 300 2340 700 2480
rect 780 2340 1100 2540
rect -210 2320 1100 2340
rect -500 2300 1100 2320
rect 1300 2560 2900 2700
rect 1300 2360 1550 2560
rect 1650 2540 2900 2560
rect 1650 2360 2040 2540
rect 1300 2340 2040 2360
rect 2120 2520 2900 2540
rect 2120 2340 2560 2520
rect 1300 2320 2560 2340
rect 2640 2320 2900 2520
rect 1300 2300 2900 2320
rect 3120 1710 3630 1810
rect -1000 1520 2600 1600
rect -1000 1500 340 1520
rect -1000 1380 -180 1500
rect -120 1380 100 1500
rect 160 1400 340 1500
rect 400 1500 2600 1520
rect 400 1400 620 1500
rect 160 1380 620 1400
rect 680 1380 2600 1500
rect -1000 1300 2600 1380
rect 3110 1036 3630 1710
rect -1000 940 2600 1000
rect -1000 920 2460 940
rect -1000 900 1940 920
rect -1000 780 1660 900
rect 1720 800 1940 900
rect 2000 800 2180 920
rect 2240 820 2460 920
rect 2520 820 2600 940
rect 2240 800 2600 820
rect 1720 780 2600 800
rect -1000 700 2600 780
rect 3110 966 3166 1036
rect 3598 966 3630 1036
rect 3110 770 3630 966
rect 5530 1636 6050 2390
rect 5530 1566 5566 1636
rect 5998 1566 6050 1636
rect 5530 1036 6050 1566
rect 5530 966 5566 1036
rect 5998 966 6050 1036
rect 3110 670 3620 770
rect 5530 750 6050 966
rect 3200 510 3500 670
rect 3120 400 3180 410
rect -600 290 2700 400
rect 2900 290 3120 400
rect -600 260 3120 290
rect -600 250 2290 260
rect -600 100 -60 250
rect 40 120 450 250
rect 560 240 2290 250
rect 560 120 1770 240
rect 40 110 1770 120
rect 1890 130 2290 240
rect 2410 130 3120 260
rect 1890 110 3120 130
rect 40 100 3120 110
rect -600 70 3120 100
rect -600 0 2700 70
rect 2900 30 3120 70
rect 3180 30 3190 400
rect 3250 300 3500 510
rect 3250 90 3260 300
rect 3320 270 4350 300
rect 3320 130 4280 270
rect 4340 130 4350 270
rect 3320 90 4350 130
rect 3120 20 3180 30
rect 3250 0 4350 90
rect 3250 -100 3500 0
use sky130_fd_pr__nfet_01v8_lvt_TV58K7  sky130_fd_pr__nfet_01v8_lvt_TV58K7_0
timestamp 1713539272
transform 1 0 2083 0 1 1410
box -683 -1810 683 1810
use sky130_fd_pr__pfet_01v8_6HGTAW  sky130_fd_pr__pfet_01v8_6HGTAW_0
timestamp 1713540189
transform 1 0 4425 0 1 7819
box -425 -1819 425 1819
use sky130_fd_pr__nfet_01v8_lvt_HS3BL4  XM1
timestamp 1713539272
transform 1 0 -104 0 1 4610
box -296 -1010 296 1010
use sky130_fd_pr__nfet_01v8_lvt_HS3BL4  XM2
timestamp 1713539272
transform 1 0 696 0 1 4610
box -296 -1010 296 1010
use sky130_fd_pr__nfet_01v8_lvt_HS3BL4  XM3
timestamp 1713539272
transform 1 0 1696 0 1 4610
box -296 -1010 296 1010
use sky130_fd_pr__nfet_01v8_lvt_HS3BL4  XM4
timestamp 1713539272
transform 1 0 2496 0 1 4610
box -296 -1010 296 1010
use sky130_fd_pr__nfet_01v8_lvt_TV58K7  XM5
timestamp 1713539272
transform 1 0 247 0 1 1448
box -683 -1810 683 1810
use sky130_fd_pr__pfet_01v8_6HGTAW  XM7
timestamp 1713540189
transform 1 0 2025 0 1 7819
box -425 -1819 425 1819
use sky130_fd_pr__pfet_01v8_3H68VM  XM8
timestamp 1713539272
transform 1 0 -22 0 1 6669
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_3H68VM  XM9
timestamp 1713539272
transform 1 0 896 0 1 6655
box -296 -619 296 619
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM10
timestamp 1713539272
transform 1 0 3296 0 1 210
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM11
timestamp 1713539272
transform 1 0 4296 0 1 210
box -296 -410 296 410
use sky130_fd_pr__pfet_01v8_6HGTAW  XM12
timestamp 1713540189
transform 1 0 3225 0 1 7819
box -425 -1819 425 1819
use sky130_fd_pr__nfet_01v8_lvt_XA7BLB  XM13
timestamp 1713540189
transform 1 0 4425 0 1 3810
box -425 -1810 425 1810
use sky130_fd_pr__nfet_01v8_lvt_7WXQKD  XM14
timestamp 1713539272
transform 1 0 3496 0 1 3810
box -296 -1810 296 1810
use sky130_fd_pr__res_xhigh_po_0p35_KNBXRF  XR1
timestamp 1713539272
transform 0 -1 4582 1 0 1601
box -201 -1582 201 1582
use sky130_fd_pr__res_xhigh_po_0p35_KNBXRF  XR4
timestamp 1713539272
transform 0 -1 4582 1 0 1001
box -201 -1582 201 1582
<< labels >>
flabel metal2 -1000 700 -680 1000 0 FreeSans 1600 0 0 0 VRF_N
port 3 nsew
flabel metal2 -1000 1300 -680 1600 0 FreeSans 1600 0 0 0 VRF
port 2 nsew
flabel metal2 -1000 4600 -800 4800 0 FreeSans 1600 0 0 0 VLO
port 0 nsew
flabel metal2 -1000 4300 -800 4500 0 FreeSans 1600 0 0 0 VLO_N
port 1 nsew
flabel metal2 -1000 4900 -800 5100 0 FreeSans 1600 0 0 0 VOUT_P
flabel metal2 -1000 5200 -800 5400 0 FreeSans 1600 0 0 0 VOUT
<< end >>
