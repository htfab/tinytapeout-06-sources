magic
tech sky130A
timestamp 1713387278
<< end >>
