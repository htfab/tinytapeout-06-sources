magic
tech sky130A
timestamp 1713041211
<< nwell >>
rect -341 -192 341 192
<< pmos >>
rect -243 -82 -143 118
rect -114 -82 -14 118
rect 14 -82 114 118
rect 143 -82 243 118
<< pdiff >>
rect -272 112 -243 118
rect -272 -76 -266 112
rect -249 -76 -243 112
rect -272 -82 -243 -76
rect -143 112 -114 118
rect -143 -76 -137 112
rect -120 -76 -114 112
rect -143 -82 -114 -76
rect -14 112 14 118
rect -14 -76 -8 112
rect 8 -76 14 112
rect -14 -82 14 -76
rect 114 112 143 118
rect 114 -76 120 112
rect 137 -76 143 112
rect 114 -82 143 -76
rect 243 112 272 118
rect 243 -76 249 112
rect 266 -76 272 112
rect 243 -82 272 -76
<< pdiffc >>
rect -266 -76 -249 112
rect -137 -76 -120 112
rect -8 -76 8 112
rect 120 -76 137 112
rect 249 -76 266 112
<< nsubdiff >>
rect -323 157 -275 174
rect 275 157 323 174
rect -323 125 -306 157
rect -323 -157 -306 -125
rect 306 -157 323 157
rect -323 -174 323 -157
<< nsubdiffcont >>
rect -275 157 275 174
rect -323 -125 -306 125
<< poly >>
rect -243 118 -143 131
rect -114 118 -14 131
rect 14 118 114 131
rect 143 118 243 131
rect -243 -105 -143 -82
rect -243 -122 -235 -105
rect -151 -122 -143 -105
rect -243 -130 -143 -122
rect -114 -105 -14 -82
rect -114 -122 -106 -105
rect -22 -122 -14 -105
rect -114 -130 -14 -122
rect 14 -105 114 -82
rect 14 -122 22 -105
rect 106 -122 114 -105
rect 14 -130 114 -122
rect 143 -105 243 -82
rect 143 -122 151 -105
rect 235 -122 243 -105
rect 143 -130 243 -122
<< polycont >>
rect -235 -122 -151 -105
rect -106 -122 -22 -105
rect 22 -122 106 -105
rect 151 -122 235 -105
<< locali >>
rect -323 157 -275 174
rect 275 157 323 174
rect -266 112 -249 120
rect -266 -84 -249 -76
rect -137 112 -120 120
rect -137 -84 -120 -76
rect -8 112 8 120
rect -8 -84 8 -76
rect 120 112 137 120
rect 120 -84 137 -76
rect 249 112 266 120
rect 249 -84 266 -76
rect -243 -122 -235 -105
rect -151 -122 -143 -105
rect -114 -122 -106 -105
rect -22 -122 -14 -105
rect 14 -122 22 -105
rect 106 -122 114 -105
rect 143 -122 151 -105
rect 235 -122 243 -105
rect 306 -157 323 157
rect -323 -174 323 -157
<< viali >>
rect -323 125 -306 157
rect -323 -125 -306 125
rect -266 28 -249 103
rect -137 -67 -120 7
rect -8 28 8 103
rect 120 -67 137 7
rect 249 28 266 103
rect -235 -122 -151 -105
rect -106 -122 -22 -105
rect 22 -122 106 -105
rect 151 -122 235 -105
rect -323 -157 -306 -125
<< metal1 >>
rect -326 157 -303 163
rect -326 -157 -323 157
rect -306 -157 -303 157
rect -269 103 -246 109
rect -269 28 -266 103
rect -249 28 -246 103
rect -269 22 -246 28
rect -11 103 11 109
rect -11 28 -8 103
rect 8 28 11 103
rect -11 22 11 28
rect 246 103 269 109
rect 246 28 249 103
rect 266 28 269 103
rect 246 22 269 28
rect -140 7 -117 13
rect -140 -67 -137 7
rect -120 -67 -117 7
rect -140 -73 -117 -67
rect 117 7 140 13
rect 117 -67 120 7
rect 137 -67 140 7
rect 117 -73 140 -67
rect -241 -105 -145 -102
rect -241 -122 -235 -105
rect -151 -122 -145 -105
rect -241 -125 -145 -122
rect -112 -105 -16 -102
rect -112 -122 -106 -105
rect -22 -122 -16 -105
rect -112 -125 -16 -122
rect 16 -105 112 -102
rect 16 -122 22 -105
rect 106 -122 112 -105
rect 16 -125 112 -122
rect 145 -105 241 -102
rect 145 -122 151 -105
rect 235 -122 241 -105
rect 145 -125 241 -122
rect -326 -163 -303 -157
<< properties >>
string FIXED_BBOX -315 -165 315 165
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 100 viagt 0
<< end >>
