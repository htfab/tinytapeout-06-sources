magic
tech sky130A
magscale 1 2
timestamp 1713540189
<< pwell >>
rect -425 -1810 425 1810
<< nmoslvt >>
rect -229 -1600 -29 1600
rect 29 -1600 229 1600
<< ndiff >>
rect -287 1588 -229 1600
rect -287 -1588 -275 1588
rect -241 -1588 -229 1588
rect -287 -1600 -229 -1588
rect -29 1588 29 1600
rect -29 -1588 -17 1588
rect 17 -1588 29 1588
rect -29 -1600 29 -1588
rect 229 1588 287 1600
rect 229 -1588 241 1588
rect 275 -1588 287 1588
rect 229 -1600 287 -1588
<< ndiffc >>
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
<< psubdiff >>
rect -389 1740 -293 1774
rect 293 1740 389 1774
rect -389 1678 -355 1740
rect 355 1678 389 1740
rect -389 -1740 -355 -1678
rect 355 -1740 389 -1678
rect -389 -1774 -293 -1740
rect 293 -1774 389 -1740
<< psubdiffcont >>
rect -293 1740 293 1774
rect -389 -1678 -355 1678
rect 355 -1678 389 1678
rect -293 -1774 293 -1740
<< poly >>
rect -229 1672 -29 1688
rect -229 1638 -213 1672
rect -45 1638 -29 1672
rect -229 1600 -29 1638
rect 29 1672 229 1688
rect 29 1638 45 1672
rect 213 1638 229 1672
rect 29 1600 229 1638
rect -229 -1638 -29 -1600
rect -229 -1672 -213 -1638
rect -45 -1672 -29 -1638
rect -229 -1688 -29 -1672
rect 29 -1638 229 -1600
rect 29 -1672 45 -1638
rect 213 -1672 229 -1638
rect 29 -1688 229 -1672
<< polycont >>
rect -213 1638 -45 1672
rect 45 1638 213 1672
rect -213 -1672 -45 -1638
rect 45 -1672 213 -1638
<< locali >>
rect -389 1740 -293 1774
rect 293 1740 389 1774
rect -389 1678 -355 1740
rect 355 1678 389 1740
rect -229 1638 -213 1672
rect -45 1638 -29 1672
rect 29 1638 45 1672
rect 213 1638 229 1672
rect -275 1588 -241 1604
rect -275 -1604 -241 -1588
rect -17 1588 17 1604
rect -17 -1604 17 -1588
rect 241 1588 275 1604
rect 241 -1604 275 -1588
rect -229 -1672 -213 -1638
rect -45 -1672 -29 -1638
rect 29 -1672 45 -1638
rect 213 -1672 229 -1638
rect -389 -1740 -355 -1678
rect 355 -1740 389 -1678
rect -389 -1774 -293 -1740
rect 293 -1774 389 -1740
<< viali >>
rect -213 1638 -45 1672
rect 45 1638 213 1672
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
rect -213 -1672 -45 -1638
rect 45 -1672 213 -1638
<< metal1 >>
rect -225 1672 -33 1678
rect -225 1638 -213 1672
rect -45 1638 -33 1672
rect -225 1632 -33 1638
rect 33 1672 225 1678
rect 33 1638 45 1672
rect 213 1638 225 1672
rect 33 1632 225 1638
rect -281 1588 -235 1600
rect -281 -1588 -275 1588
rect -241 -1588 -235 1588
rect -281 -1600 -235 -1588
rect -23 1588 23 1600
rect -23 -1588 -17 1588
rect 17 -1588 23 1588
rect -23 -1600 23 -1588
rect 235 1588 281 1600
rect 235 -1588 241 1588
rect 275 -1588 281 1588
rect 235 -1600 281 -1588
rect -225 -1638 -33 -1632
rect -225 -1672 -213 -1638
rect -45 -1672 -33 -1638
rect -225 -1678 -33 -1672
rect 33 -1638 225 -1632
rect 33 -1672 45 -1638
rect 213 -1672 225 -1638
rect 33 -1678 225 -1672
<< properties >>
string FIXED_BBOX -372 -1757 372 1757
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 16.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
