* NGSPICE file created from vbias_resistor_parax.ext - technology: sky130A

.subckt vbias_resistor_parax VDD VSS VBIAS
X0 VDD VBIAS VSS.t8 sky130_fd_pr__res_xhigh_po_0p35 l=2.8
X1 VBIAS.t3 VBIAS.t2 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X2 VSS.t5 VBIAS.t0 VBIAS.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X3 VSS.t3 VBIAS.t4 VBIAS.t5 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X4 VBIAS.t7 VBIAS.t6 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
R0 VBIAS.n1 VBIAS.n0 66.318
R1 VBIAS.n4 VBIAS.n3 66.3172
R2 VBIAS.n4 VBIAS.t2 25.5777
R3 VBIAS.n5 VBIAS.t4 25.5624
R4 VBIAS.n1 VBIAS.t6 25.5552
R5 VBIAS.n2 VBIAS.t0 25.5479
R6 VBIAS.n3 VBIAS.t5 17.4005
R7 VBIAS.n3 VBIAS.t3 17.4005
R8 VBIAS.n0 VBIAS.t1 17.4005
R9 VBIAS.n0 VBIAS.t7 17.4005
R10 VBIAS VBIAS.n6 0.550632
R11 VBIAS.n6 VBIAS.n2 0.247722
R12 VBIAS.n6 VBIAS.n5 0.205547
R13 VBIAS.n2 VBIAS.n1 0.00582231
R14 VBIAS.n5 VBIAS.n4 0.00162952
R15 VSS.n19 VSS.n8 7358.53
R16 VSS.n21 VSS.n8 7358.53
R17 VSS.n21 VSS.n7 7358.53
R18 VSS.n19 VSS.n7 7358.53
R19 VSS.n16 VSS.n15 5446.47
R20 VSS.n16 VSS.n11 5446.47
R21 VSS.n14 VSS.n11 5446.47
R22 VSS.n15 VSS.n14 5446.47
R23 VSS.t6 VSS.t2 569.909
R24 VSS.t4 VSS.t0 569.909
R25 VSS.t2 VSS.n7 543.811
R26 VSS.t0 VSS.n8 543.811
R27 VSS.n18 VSS.n11 301.05
R28 VSS.n15 VSS.n12 292.5
R29 VSS.n15 VSS.t8 292.5
R30 VSS.n11 VSS.t8 292.5
R31 VSS.n13 VSS.t8 184.163
R32 VSS.n9 VSS.t4 150.566
R33 VSS.n20 VSS.n9 134.389
R34 VSS.n7 VSS.n5 117.001
R35 VSS.n8 VSS.n6 117.001
R36 VSS.n3 VSS.t1 85.0617
R37 VSS.n0 VSS.t3 85.0584
R38 VSS.n2 VSS.n1 67.1938
R39 VSS.n17 VSS.n12 58.9599
R40 VSS.n12 VSS.n10 58.8533
R41 VSS.n13 VSS.t6 51.0186
R42 VSS.n20 VSS.t8 49.7743
R43 VSS.n22 VSS.n6 41.3952
R44 VSS.n23 VSS.n5 33.8916
R45 VSS.n19 VSS.n18 29.443
R46 VSS.n14 VSS.n10 27.8576
R47 VSS.n14 VSS.n13 27.8576
R48 VSS.n17 VSS.n16 27.8576
R49 VSS.n16 VSS.n9 27.8576
R50 VSS.n18 VSS.n6 22.4993
R51 VSS.n20 VSS.n19 20.8934
R52 VSS.n22 VSS.n21 20.8934
R53 VSS.n21 VSS.n20 20.8934
R54 VSS.n1 VSS.t7 17.4005
R55 VSS.n1 VSS.t5 17.4005
R56 VSS.n18 VSS.n5 14.8536
R57 VSS.n18 VSS.n17 11.7279
R58 VSS.n18 VSS.n10 11.5983
R59 VSS.n4 VSS.n0 4.50515
R60 VSS.n23 VSS.n22 0.778615
R61 VSS.n4 VSS.n3 0.0780862
R62 VSS.n24 VSS.n23 0.0646379
R63 VSS VSS.n24 0.0151861
R64 VSS.n24 VSS.n4 0.00548879
R65 VSS.n2 VSS.n0 0.00251613
R66 VSS.n3 VSS.n2 0.00150806
C0 VBIAS VDD 0.049588f
.ends

