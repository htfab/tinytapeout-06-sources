magic
tech sky130A
magscale 1 2
timestamp 1713057736
<< nwell >>
rect -425 -1231 425 1231
<< pmos >>
rect -229 683 -29 1083
rect 29 683 229 1083
rect -229 118 -29 518
rect 29 118 229 518
rect -229 -447 -29 -47
rect 29 -447 229 -47
rect -229 -1012 -29 -612
rect 29 -1012 229 -612
<< pdiff >>
rect -287 1071 -229 1083
rect -287 695 -275 1071
rect -241 695 -229 1071
rect -287 683 -229 695
rect -29 1071 29 1083
rect -29 695 -17 1071
rect 17 695 29 1071
rect -29 683 29 695
rect 229 1071 287 1083
rect 229 695 241 1071
rect 275 695 287 1071
rect 229 683 287 695
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect -287 -59 -229 -47
rect -287 -435 -275 -59
rect -241 -435 -229 -59
rect -287 -447 -229 -435
rect -29 -59 29 -47
rect -29 -435 -17 -59
rect 17 -435 29 -59
rect -29 -447 29 -435
rect 229 -59 287 -47
rect 229 -435 241 -59
rect 275 -435 287 -59
rect 229 -447 287 -435
rect -287 -624 -229 -612
rect -287 -1000 -275 -624
rect -241 -1000 -229 -624
rect -287 -1012 -229 -1000
rect -29 -624 29 -612
rect -29 -1000 -17 -624
rect 17 -1000 29 -624
rect -29 -1012 29 -1000
rect 229 -624 287 -612
rect 229 -1000 241 -624
rect 275 -1000 287 -624
rect 229 -1012 287 -1000
<< pdiffc >>
rect -275 695 -241 1071
rect -17 695 17 1071
rect 241 695 275 1071
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect -275 -1000 -241 -624
rect -17 -1000 17 -624
rect 241 -1000 275 -624
<< nsubdiff >>
rect -389 1161 -293 1195
rect 293 1161 389 1195
rect -389 -1161 -355 1161
rect 355 -1161 389 1161
rect -389 -1195 389 -1161
<< nsubdiffcont >>
rect -293 1161 293 1195
<< poly >>
rect -229 1083 -29 1109
rect 29 1083 229 1109
rect -229 636 -29 683
rect -229 602 -213 636
rect -45 602 -29 636
rect -229 586 -29 602
rect 29 636 229 683
rect 29 602 45 636
rect 213 602 229 636
rect 29 586 229 602
rect -229 518 -29 544
rect 29 518 229 544
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -47 -29 -21
rect 29 -47 229 -21
rect -229 -494 -29 -447
rect -229 -528 -213 -494
rect -45 -528 -29 -494
rect -229 -544 -29 -528
rect 29 -494 229 -447
rect 29 -528 45 -494
rect 213 -528 229 -494
rect 29 -544 229 -528
rect -229 -612 -29 -586
rect 29 -612 229 -586
rect -229 -1059 -29 -1012
rect -229 -1093 -213 -1059
rect -45 -1093 -29 -1059
rect -229 -1109 -29 -1093
rect 29 -1059 229 -1012
rect 29 -1093 45 -1059
rect 213 -1093 229 -1059
rect 29 -1109 229 -1093
<< polycont >>
rect -213 602 -45 636
rect 45 602 213 636
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -528 -45 -494
rect 45 -528 213 -494
rect -213 -1093 -45 -1059
rect 45 -1093 213 -1059
<< locali >>
rect -389 -1161 -355 1195
rect -275 1071 -241 1087
rect -275 679 -241 695
rect -17 1071 17 1087
rect -17 679 17 695
rect 241 1071 275 1087
rect 241 679 275 695
rect -229 602 -213 636
rect -45 602 -29 636
rect 29 602 45 636
rect 213 602 229 636
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -275 -59 -241 -43
rect -275 -451 -241 -435
rect -17 -59 17 -43
rect -17 -451 17 -435
rect 241 -59 275 -43
rect 241 -451 275 -435
rect -229 -528 -213 -494
rect -45 -528 -29 -494
rect 29 -528 45 -494
rect 213 -528 229 -494
rect -275 -624 -241 -608
rect -275 -1016 -241 -1000
rect -17 -624 17 -608
rect -17 -1016 17 -1000
rect 241 -624 275 -608
rect 241 -1016 275 -1000
rect -229 -1093 -213 -1059
rect -45 -1093 -29 -1059
rect 29 -1093 45 -1059
rect 213 -1093 229 -1059
rect 355 -1161 389 1195
rect -389 -1195 389 -1161
<< viali >>
rect -355 1161 -293 1195
rect -293 1161 293 1195
rect 293 1161 355 1195
rect -275 695 -241 1071
rect -17 695 17 1071
rect 241 695 275 1071
rect -213 602 -45 636
rect 45 602 213 636
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -213 37 -45 71
rect 45 37 213 71
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect -213 -528 -45 -494
rect 45 -528 213 -494
rect -275 -1000 -241 -624
rect -17 -1000 17 -624
rect 241 -1000 275 -624
rect -213 -1093 -45 -1059
rect 45 -1093 213 -1059
<< metal1 >>
rect -367 1195 367 1201
rect -367 1161 -355 1195
rect 355 1161 367 1195
rect -367 1155 367 1161
rect -281 1071 -235 1083
rect -281 695 -275 1071
rect -241 695 -235 1071
rect -281 683 -235 695
rect -23 1071 23 1083
rect -23 695 -17 1071
rect 17 695 23 1071
rect -23 683 23 695
rect 235 1071 281 1083
rect 235 695 241 1071
rect 275 695 281 1071
rect 235 683 281 695
rect -225 636 -33 642
rect -225 602 -213 636
rect -45 602 -33 636
rect -225 596 -33 602
rect 33 636 225 642
rect 33 602 45 636
rect 213 602 225 636
rect 33 596 225 602
rect -281 506 -235 518
rect -281 130 -275 506
rect -241 130 -235 506
rect -281 118 -235 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 235 506 281 518
rect 235 130 241 506
rect 275 130 281 506
rect 235 118 281 130
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -281 -59 -235 -47
rect -281 -435 -275 -59
rect -241 -435 -235 -59
rect -281 -447 -235 -435
rect -23 -59 23 -47
rect -23 -435 -17 -59
rect 17 -435 23 -59
rect -23 -447 23 -435
rect 235 -59 281 -47
rect 235 -435 241 -59
rect 275 -435 281 -59
rect 235 -447 281 -435
rect -225 -494 -33 -488
rect -225 -528 -213 -494
rect -45 -528 -33 -494
rect -225 -534 -33 -528
rect 33 -494 225 -488
rect 33 -528 45 -494
rect 213 -528 225 -494
rect 33 -534 225 -528
rect -281 -624 -235 -612
rect -281 -1000 -275 -624
rect -241 -1000 -235 -624
rect -281 -1012 -235 -1000
rect -23 -624 23 -612
rect -23 -1000 -17 -624
rect 17 -1000 23 -624
rect -23 -1012 23 -1000
rect 235 -624 281 -612
rect 235 -1000 241 -624
rect 275 -1000 281 -624
rect 235 -1012 281 -1000
rect -225 -1059 -33 -1053
rect -225 -1093 -213 -1059
rect -45 -1093 -33 -1059
rect -225 -1099 -33 -1093
rect 33 -1059 225 -1053
rect 33 -1093 45 -1059
rect 213 -1093 225 -1059
rect 33 -1099 225 -1093
<< properties >>
string FIXED_BBOX -372 -1178 372 1178
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 2 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
