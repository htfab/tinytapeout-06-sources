magic
tech sky130A
magscale 1 2
timestamp 1713432866
<< error_p >>
rect -31 531 31 537
rect -31 497 -19 531
rect -31 491 31 497
rect -31 -497 31 -491
rect -31 -531 -19 -497
rect -31 -537 31 -531
<< nwell >>
rect -231 -669 231 669
<< pmoslvt >>
rect -35 -450 35 450
<< pdiff >>
rect -93 438 -35 450
rect -93 -438 -81 438
rect -47 -438 -35 438
rect -93 -450 -35 -438
rect 35 438 93 450
rect 35 -438 47 438
rect 81 -438 93 438
rect 35 -450 93 -438
<< pdiffc >>
rect -81 -438 -47 438
rect 47 -438 81 438
<< nsubdiff >>
rect -195 599 -99 633
rect 99 599 195 633
rect -195 537 -161 599
rect 161 537 195 599
rect -195 -599 -161 -537
rect 161 -599 195 -537
rect -195 -633 -99 -599
rect 99 -633 195 -599
<< nsubdiffcont >>
rect -99 599 99 633
rect -195 -537 -161 537
rect 161 -537 195 537
rect -99 -633 99 -599
<< poly >>
rect -35 531 35 547
rect -35 497 -19 531
rect 19 497 35 531
rect -35 450 35 497
rect -35 -497 35 -450
rect -35 -531 -19 -497
rect 19 -531 35 -497
rect -35 -547 35 -531
<< polycont >>
rect -19 497 19 531
rect -19 -531 19 -497
<< locali >>
rect -195 599 -99 633
rect 99 599 195 633
rect -195 537 -161 599
rect 161 537 195 599
rect -35 497 -19 531
rect 19 497 35 531
rect -81 438 -47 454
rect -81 -454 -47 -438
rect 47 438 81 454
rect 47 -454 81 -438
rect -35 -531 -19 -497
rect 19 -531 35 -497
rect -195 -599 -161 -537
rect 161 -599 195 -537
rect -195 -633 -99 -599
rect 99 -633 195 -599
<< viali >>
rect -19 497 19 531
rect -81 -438 -47 438
rect 47 -438 81 438
rect -19 -531 19 -497
<< metal1 >>
rect -31 531 31 537
rect -31 497 -19 531
rect 19 497 31 531
rect -31 491 31 497
rect -87 438 -41 450
rect -87 -438 -81 438
rect -47 -438 -41 438
rect -87 -450 -41 -438
rect 41 438 87 450
rect 41 -438 47 438
rect 81 -438 87 438
rect 41 -450 87 -438
rect -31 -497 31 -491
rect -31 -531 -19 -497
rect 19 -531 31 -497
rect -31 -537 31 -531
<< properties >>
string FIXED_BBOX -178 -616 178 616
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4.5 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
