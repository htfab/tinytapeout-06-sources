** sch_path: /foss/designs/flash-adc/xschem/adc_with_encoder.sch
.subckt adc_with_encoder VDD OUT3 OUT2 IN OUT1 OUT0 VSS
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT0
*.opin OUT1
*.opin OUT2
*.opin OUT3
x1 VDD IN net1 net2 net3 net4 net5 net6 net7 net8 net9 net10 net11 net12 net13 net14 net15 VSS flash_adc
x2 net1 VDD net2 net3 net4 net5 net6 net7 net8 OUT3 net9 OUT2 net10 OUT1 net11 OUT0 net12 net13 net14 VSS net15 encoder_tree
.ends

* expanding   symbol:  /foss/designs/flash-adc/xschem/flash_adc.sym # of pins=18
** sym_path: /foss/designs/flash-adc/xschem/flash_adc.sym
** sch_path: /foss/designs/flash-adc/xschem/flash_adc.sch
.subckt flash_adc VDD IN OUT14 OUT13 OUT12 OUT11 OUT10 OUT9 OUT8 OUT7 OUT6 OUT5 OUT4 OUT3 OUT2 OUT1 OUT0 VSS
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT0
*.opin OUT1
*.opin OUT2
*.opin OUT3
*.opin OUT4
*.opin OUT5
*.opin OUT6
*.opin OUT7
*.opin OUT8
*.opin OUT9
*.opin OUT10
*.opin OUT11
*.opin OUT12
*.opin OUT13
*.opin OUT14
x1 VDD net2 IN VSS vfollower
x2 VDD net1 IN VSS vfollower
x3 VDD net3 IN VSS vfollower
x4 VDD net4 IN VSS vfollower
x5 net10 VDD net2 OUT0 VSS VSS ladder_rung
x6 net9 VDD net2 OUT1 VSS net10 ladder_rung
x7 net8 VDD net2 OUT2 VSS net9 ladder_rung
x8 net5 VDD net2 OUT3 VSS net8 ladder_rung
x9 net13 VDD net1 OUT4 VSS net5 ladder_rung
x10 net12 VDD net1 OUT5 VSS net13 ladder_rung
x11 net11 VDD net1 OUT6 VSS net12 ladder_rung
x12 net6 VDD net1 OUT7 VSS net11 ladder_rung
x13 net16 VDD net3 OUT8 VSS net6 ladder_rung
x14 net15 VDD net3 OUT9 VSS net16 ladder_rung
x15 net14 VDD net3 OUT10 VSS net15 ladder_rung
x16 net7 VDD net3 OUT11 VSS net14 ladder_rung
x17 net18 VDD net4 OUT12 VSS net7 ladder_rung
x18 net17 VDD net4 OUT13 VSS net18 ladder_rung
x19 VDD VDD net4 OUT14 VSS net17 ladder_rung
.ends


* expanding   symbol:  /foss/designs/flash-adc/xschem/encoder_tree.sym # of pins=21
** sym_path: /foss/designs/flash-adc/xschem/encoder_tree.sym
** sch_path: /foss/designs/flash-adc/xschem/encoder_tree.sch
.subckt encoder_tree IN14 VDD IN13 IN12 IN11 IN10 IN9 IN8 IN7 OUT3 IN6 OUT2 IN5 OUT1 IN4 OUT0 IN3 IN2 IN1 VSS IN0
*.ipin IN0
*.ipin IN1
*.ipin IN2
*.ipin IN3
*.ipin IN4
*.ipin IN5
*.ipin IN6
*.ipin IN7
*.ipin IN8
*.ipin IN9
*.ipin IN10
*.ipin IN11
*.ipin IN12
*.ipin IN13
*.ipin IN14
*.opin OUT0
*.opin OUT1
*.opin OUT2
*.opin OUT3
*.iopin VDD
*.iopin VSS
x1 IN2 IN1 IN0 VSS VSS VDD VDD net3 sky130_fd_sc_hd__maj3_4
x2 IN4 IN3 IN2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__maj3_4
x3 IN6 IN5 IN4 VSS VSS VDD VDD net4 sky130_fd_sc_hd__maj3_4
x4 IN8 IN7 IN6 VSS VSS VDD VDD net8 sky130_fd_sc_hd__maj3_4
x5 IN10 IN9 IN8 VSS VSS VDD VDD net9 sky130_fd_sc_hd__maj3_4
x6 IN12 IN11 IN10 VSS VSS VDD VDD net11 sky130_fd_sc_hd__maj3_4
x7 IN14 IN13 IN12 VSS VSS VDD VDD net10 sky130_fd_sc_hd__maj3_4
x8 IN0 IN2 net3 VSS VSS VDD VDD net7 sky130_fd_sc_hd__mux2_4
x9 IN4 IN6 net4 VSS VSS VDD VDD net6 sky130_fd_sc_hd__mux2_4
x10 IN8 IN10 net9 VSS VSS VDD VDD net13 sky130_fd_sc_hd__mux2_4
x11 IN12 IN14 net10 VSS VSS VDD VDD net14 sky130_fd_sc_hd__mux2_4
x12 net4 net1 net3 VSS VSS VDD VDD net2 sky130_fd_sc_hd__maj3_4
x13 net9 net8 net4 VSS VSS VDD VDD net15 sky130_fd_sc_hd__maj3_4
x14 net10 net11 net9 VSS VSS VDD VDD net12 sky130_fd_sc_hd__maj3_4
x15 net3 net4 net2 VSS VSS VDD VDD net5 sky130_fd_sc_hd__mux2_4
x16 net7 net6 net2 VSS VSS VDD VDD net18 sky130_fd_sc_hd__mux2_4
x17 net9 net10 net12 VSS VSS VDD VDD net16 sky130_fd_sc_hd__mux2_4
x18 net13 net14 net12 VSS VSS VDD VDD net17 sky130_fd_sc_hd__mux2_4
x19 net12 net15 net2 VSS VSS VDD VDD OUT3 sky130_fd_sc_hd__maj3_4
x20 net2 net12 OUT3 VSS VSS VDD VDD OUT2 sky130_fd_sc_hd__mux2_4
x21 net5 net16 OUT3 VSS VSS VDD VDD OUT1 sky130_fd_sc_hd__mux2_4
x22 net18 net17 OUT3 VSS VSS VDD VDD OUT0 sky130_fd_sc_hd__mux2_4
.ends


* expanding   symbol:  /foss/designs/flash-adc/xschem/vfollower.sym # of pins=4
** sym_path: /foss/designs/flash-adc/xschem/vfollower.sym
** sch_path: /foss/designs/flash-adc/xschem/vfollower.sch
.subckt vfollower VDD OUT IN VSS
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
x1 VDD OUT IN OUT VSS opamp
.ends


* expanding   symbol:  /foss/designs/flash-adc/xschem/ladder_rung.sym # of pins=6
** sym_path: /foss/designs/flash-adc/xschem/ladder_rung.sym
** sch_path: /foss/designs/flash-adc/xschem/ladder_rung.sch
.subckt ladder_rung HI VDD IN OUT VSS LO
*.opin OUT
*.iopin VDD
*.iopin VSS
*.ipin IN
*.iopin LO
*.iopin HI
XR1 LO net1 VSS sky130_fd_pr__res_xhigh_po_0p35 L=2.34 mult=1 m=1
x5 VDD OUT IN net1 VSS comparator
XR2 net1 HI VSS sky130_fd_pr__res_xhigh_po_0p35 L=2.34 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/flash-adc/xschem/opamp.sym # of pins=5
** sym_path: /foss/designs/flash-adc/xschem/opamp.sym
** sch_path: /foss/designs/flash-adc/xschem/opamp.sch
.subckt opamp VDD OUT P N VSS
*.iopin VDD
*.iopin VSS
*.ipin P
*.ipin N
*.opin OUT
XR1 net2 VDD VSS sky130_fd_pr__res_xhigh_po_0p35 L=24.36 mult=1 m=1
XM1 net2 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM7 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM8 OUT net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM4 net6 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 net1 P net6 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM6 OUT N net6 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 net5 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM9 net4 net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 VDD net5 net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM10 net3 P net4 VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM11 OUT N net4 VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM12 net3 net3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM13 OUT net3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  /foss/designs/flash-adc/xschem/comparator.sym # of pins=5
** sym_path: /foss/designs/flash-adc/xschem/comparator.sym
** sch_path: /foss/designs/flash-adc/xschem/comparator.sch
.subckt comparator VDD OUT P N VSS
*.iopin VDD
*.iopin VSS
*.ipin P
*.ipin N
*.opin OUT
x1 VDD net1 P N VSS opamp
x2 VDD OUT net1 VSS buffer
.ends


* expanding   symbol:  /foss/designs/flash-adc/xschem/buffer.sym # of pins=4
** sym_path: /foss/designs/flash-adc/xschem/buffer.sym
** sch_path: /foss/designs/flash-adc/xschem/buffer.sch
.subckt buffer VDD OUT IN VSS
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 net1 IN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 IN VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
