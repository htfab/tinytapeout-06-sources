magic
tech sky130A
magscale 1 2
timestamp 1713125316
<< pwell >>
rect -468 -1372 32 -1262
rect -962 -2040 -586 -1898
<< locali >>
rect -1652 -136 -1470 -122
rect -1652 -192 -1638 -136
rect -1482 -192 -1470 -136
rect -1652 -924 -1470 -192
rect -1652 -1062 -1468 -924
rect -1650 -1260 -1470 -1062
rect -1650 -1380 -1614 -1260
rect -1504 -1380 -1470 -1260
rect -1650 -1420 -1470 -1380
<< viali >>
rect -418 140 -14 174
rect 1134 140 1520 174
rect 3406 10 3604 44
rect -1638 -192 -1482 -136
rect -420 -642 -14 -608
rect 1264 -642 1440 -608
rect -1614 -1380 -1504 -1260
rect 2394 -1358 2488 -1324
rect -356 -1564 -46 -1530
rect 1250 -1564 1460 -1530
rect 3224 -1822 3736 -1788
rect -900 -1950 -648 -1916
rect -2028 -3364 -1776 -3330
<< metal1 >>
rect -2676 584 3844 600
rect -2676 246 -2660 584
rect -2414 246 3844 584
rect -2676 224 3844 246
rect -782 174 404 224
rect -782 140 -418 174
rect -14 140 404 174
rect -782 20 404 140
rect 746 216 1940 224
rect 746 174 1938 216
rect 746 140 1134 174
rect 1520 140 1938 174
rect 746 20 1938 140
rect 1990 -8 2356 -2
rect 1990 -20 2222 -8
rect 1982 -22 2222 -20
rect -1392 -28 2222 -22
rect -1392 -98 -1384 -28
rect -1238 -64 2222 -28
rect -1238 -98 -1230 -64
rect 1990 -80 2222 -64
rect 2348 -80 2356 -8
rect 1990 -90 2356 -80
rect -1392 -106 -1230 -98
rect -1652 -134 -1470 -122
rect -788 -134 400 -114
rect -1652 -136 400 -134
rect -1652 -192 -1638 -136
rect -1482 -184 400 -136
rect -1482 -192 -1470 -184
rect -1652 -208 -1470 -192
rect -2332 -352 -2132 -284
rect 834 -324 1036 -316
rect 834 -352 846 -324
rect -2332 -420 846 -352
rect -2332 -484 -2132 -420
rect 834 -464 846 -420
rect 1026 -464 1036 -324
rect 834 -474 1036 -464
rect 1234 -508 1478 -118
rect 1858 -322 2030 -314
rect 1858 -462 1868 -322
rect 2020 -360 2030 -322
rect 2022 -414 2030 -360
rect 2020 -462 2030 -414
rect 1858 -474 2030 -462
rect -468 -572 1478 -508
rect -468 -608 28 -572
rect -468 -642 -420 -608
rect -14 -642 28 -608
rect -2328 -790 -856 -722
rect -468 -758 28 -642
rect 1234 -608 1478 -572
rect 1234 -642 1264 -608
rect 1440 -642 1478 -608
rect 1234 -754 1478 -642
rect -2328 -866 492 -790
rect 1988 -810 2028 -474
rect 662 -852 2028 -810
rect -2328 -922 -856 -866
rect 1988 -888 2028 -852
rect -2330 -1260 -1470 -1220
rect -2330 -1380 -1614 -1260
rect -1504 -1380 -1470 -1260
rect -468 -1324 32 -900
rect 1232 -1048 1480 -902
rect 2392 -944 2486 224
rect 3148 160 3844 224
rect 2922 44 4098 160
rect 2922 10 3406 44
rect 3604 10 4098 44
rect 2518 -12 2650 -6
rect 2518 -82 2526 -12
rect 2642 -82 2650 -12
rect 2518 -92 2650 -82
rect 2548 -132 2650 -92
rect 2922 -106 4098 10
rect 2548 -154 2862 -132
rect 2548 -168 3082 -154
rect 3906 -168 4188 -154
rect 2548 -200 4188 -168
rect 2548 -222 2862 -200
rect 3316 -750 3718 -248
rect 1232 -1122 2372 -1048
rect 1232 -1272 1480 -1122
rect -858 -1374 2000 -1324
rect -2330 -1420 -1470 -1380
rect -2678 -1916 -2396 -1900
rect -2678 -2248 -2660 -1916
rect -2408 -2046 -2396 -1916
rect -2408 -2124 -1812 -2046
rect -2408 -2248 -1814 -2124
rect -2678 -2260 -1814 -2248
rect -1652 -2996 -1470 -1420
rect -468 -1530 32 -1414
rect -468 -1564 -356 -1530
rect -46 -1564 32 -1530
rect -962 -1916 -586 -1898
rect -962 -1950 -900 -1916
rect -648 -1950 -586 -1916
rect -1392 -2022 -1230 -2016
rect -1392 -2026 -1382 -2022
rect -1392 -2090 -1384 -2026
rect -1236 -2038 -1230 -2022
rect -1236 -2040 -1030 -2038
rect -962 -2040 -586 -1950
rect -468 -2040 32 -1564
rect 1230 -1530 1480 -1416
rect 1230 -1564 1250 -1530
rect 1460 -1564 1480 -1530
rect 1230 -2040 1480 -1564
rect 2134 -1530 2226 -1122
rect 2418 -1258 2474 -944
rect 3316 -950 5620 -750
rect 2770 -994 3278 -978
rect 2508 -1020 2554 -1018
rect 2770 -1020 2784 -994
rect 2508 -1154 2784 -1020
rect 2770 -1208 2784 -1154
rect 3266 -1208 3278 -994
rect 2770 -1224 3278 -1208
rect 2382 -1324 2512 -1316
rect 2382 -1358 2394 -1324
rect 2488 -1358 2512 -1324
rect 2382 -1368 2512 -1358
rect 2134 -1536 2276 -1530
rect 2134 -1630 2140 -1536
rect 2268 -1630 2276 -1536
rect 2134 -1638 2276 -1630
rect 2382 -2038 2510 -1368
rect 3316 -1530 3718 -950
rect 2550 -1536 2672 -1530
rect 2550 -1632 2558 -1536
rect 2666 -1574 2672 -1536
rect 2666 -1576 2876 -1574
rect 2666 -1618 4170 -1576
rect 4970 -1612 5174 -950
rect 2666 -1632 2672 -1618
rect 2550 -1638 2672 -1632
rect 4862 -1626 5258 -1612
rect 3132 -1788 3834 -1674
rect 3132 -1822 3224 -1788
rect 3736 -1822 3834 -1788
rect 3132 -2038 3834 -1822
rect 2382 -2040 3834 -2038
rect -1392 -2094 -1382 -2090
rect -1236 -2094 3834 -2040
rect 4862 -2076 4878 -1626
rect 5238 -2076 5258 -1626
rect 4862 -2092 5258 -2076
rect -1392 -2102 3834 -2094
rect -1230 -2230 3834 -2102
rect -1230 -2552 -1030 -2230
rect -1990 -3156 -686 -2996
rect -1990 -3234 -684 -3156
rect -584 -3296 -404 -2230
rect -2160 -3330 -404 -3296
rect -2160 -3364 -2028 -3330
rect -1776 -3364 -404 -3330
rect -2160 -3472 -404 -3364
<< via1 >>
rect -2660 246 -2414 584
rect -1384 -98 -1238 -28
rect 2222 -80 2348 -8
rect 846 -464 1026 -324
rect 1868 -360 2020 -322
rect 1868 -414 2022 -360
rect 1868 -462 2020 -414
rect 2526 -82 2642 -12
rect -2660 -2248 -2408 -1916
rect -1382 -2026 -1236 -2022
rect -1384 -2090 -1236 -2026
rect 2784 -1208 3266 -994
rect 2140 -1630 2268 -1536
rect 2558 -1632 2666 -1536
rect -1382 -2094 -1236 -2090
rect 4878 -2076 5238 -1626
<< metal2 >>
rect -2676 584 -2396 600
rect -2676 246 -2660 584
rect -2414 246 -2396 584
rect -2676 -1916 -2396 246
rect 2214 -8 2356 -2
rect -2676 -2248 -2660 -1916
rect -2408 -2248 -2396 -1916
rect -1392 -28 -1230 -22
rect -1392 -98 -1384 -28
rect -1238 -98 -1230 -28
rect 2214 -80 2222 -8
rect 2348 -20 2356 -8
rect 2518 -12 2650 -6
rect 2518 -20 2526 -12
rect 2348 -64 2526 -20
rect 2348 -80 2356 -64
rect 2214 -90 2356 -80
rect 2518 -82 2526 -64
rect 2642 -82 2650 -12
rect 2518 -92 2650 -82
rect -1392 -2022 -1230 -98
rect 834 -324 1036 -316
rect 834 -464 846 -324
rect 1026 -352 1036 -324
rect 1858 -322 2030 -314
rect 1858 -352 1868 -322
rect 1026 -420 1868 -352
rect 2020 -360 2030 -322
rect 2022 -414 2030 -360
rect 1026 -464 1036 -420
rect 834 -474 1036 -464
rect 1858 -462 1868 -420
rect 2020 -462 2030 -414
rect 1858 -474 2030 -462
rect 2770 -994 3278 -978
rect 2770 -1208 2784 -994
rect 3266 -1208 3278 -994
rect 2770 -1224 3278 -1208
rect 2134 -1536 2672 -1530
rect 2134 -1630 2140 -1536
rect 2268 -1630 2558 -1536
rect 2134 -1632 2558 -1630
rect 2666 -1632 2672 -1536
rect 2134 -1638 2672 -1632
rect 4862 -1626 5258 -1612
rect -1392 -2026 -1382 -2022
rect -1392 -2090 -1384 -2026
rect -1392 -2094 -1382 -2090
rect -1236 -2094 -1230 -2022
rect 4862 -2076 4878 -1626
rect 5238 -2076 5258 -1626
rect 4862 -2092 5258 -2076
rect -1392 -2102 -1230 -2094
rect -2676 -2260 -2396 -2248
<< via2 >>
rect 2784 -1208 3266 -994
rect 4878 -2076 5238 -1626
<< metal3 >>
rect 2770 -994 3278 -978
rect 2770 -1208 2784 -994
rect 3266 -1208 3278 -994
rect 2770 -1224 3278 -1208
rect 4862 -1626 5258 -1612
rect 4862 -2076 4878 -1626
rect 5238 -2076 5258 -1626
rect 4862 -2092 5258 -2076
<< via3 >>
rect 2784 -1208 3266 -994
rect 4878 -2076 5238 -1626
<< metal4 >>
rect 2770 -994 3278 -978
rect 2770 -1208 2784 -994
rect 3266 -1022 3278 -994
rect 3266 -1156 4492 -1022
rect 3266 -1208 3278 -1156
rect 2770 -1224 3278 -1208
rect 4350 -1992 4492 -1156
rect 2736 -2140 4492 -1992
rect 4862 -1626 5258 -1612
rect 4862 -2076 4878 -1626
rect 5238 -2076 5258 -1626
rect 4862 -2092 5258 -2076
rect 2736 -2372 3104 -2140
rect 4974 -2710 5176 -2092
rect 4970 -2758 5176 -2710
rect 4970 -3584 5174 -2758
rect 3374 -4096 5176 -3584
use sky130_fd_pr__cap_mim_m3_1_QJVKAD  sky130_fd_pr__cap_mim_m3_1_QJVKAD_0
timestamp 1712676954
transform 1 0 1535 0 1 -3792
box -1941 -1540 1941 1540
use sky130_fd_pr__pfet_01v8_XPP7BA  XM1
timestamp 1712505088
transform 0 1 -189 -1 0 -828
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM2
timestamp 1712505088
transform 0 1 1343 -1 0 -828
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM3
timestamp 1712505088
transform 0 1 -186 -1 0 -1344
box -256 -810 256 810
use sky130_fd_pr__nfet_01v8_3BHWKV  XM4
timestamp 1712505088
transform 0 1 1328 -1 0 -1344
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM5
timestamp 1712505088
transform 0 1 1343 -1 0 -46
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM6
timestamp 1712505088
transform 0 1 3500 -1 0 -1602
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM7
timestamp 1712505088
transform 0 1 3509 -1 0 -176
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM8
timestamp 1712505088
transform 0 1 -189 -1 0 -46
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_7QHW3M  XM9
timestamp 1712505088
transform 1 0 2442 0 1 -1084
box -256 -310 256 310
use sky130_fd_pr__res_generic_nd_GV5DH4  XR1
timestamp 1713121488
transform 1 0 -1902 0 1 -2639
box -258 -761 258 761
use sky130_fd_pr__res_generic_nd_GV5DH4  XR2
timestamp 1713121488
transform 1 0 -774 0 1 -2641
box -258 -761 258 761
<< labels >>
flabel metal1 -1230 400 -1030 600 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -2330 -1420 -2130 -1220 0 FreeSans 256 0 0 0 ZREF
port 1 nsew
flabel metal1 -1230 -2552 -1030 -2352 0 FreeSans 256 0 0 0 VGND
port 5 nsew
flabel metal1 -2328 -922 -2128 -722 0 FreeSans 256 0 0 0 vin_n
port 2 nsew
flabel metal1 -2332 -484 -2132 -284 0 FreeSans 256 0 0 0 vin_p
port 3 nsew
flabel metal1 5420 -950 5620 -750 0 FreeSans 256 0 0 0 Vout
port 4 nsew
<< end >>
