magic
tech sky130A
magscale 1 2
timestamp 1713057736
<< nwell >>
rect -683 -666 683 666
<< pmos >>
rect -487 118 -287 518
rect -229 118 -29 518
rect 29 118 229 518
rect 287 118 487 518
rect -487 -447 -287 -47
rect -229 -447 -29 -47
rect 29 -447 229 -47
rect 287 -447 487 -47
<< pdiff >>
rect -545 506 -487 518
rect -545 130 -533 506
rect -499 130 -487 506
rect -545 118 -487 130
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect 487 506 545 518
rect 487 130 499 506
rect 533 130 545 506
rect 487 118 545 130
rect -545 -59 -487 -47
rect -545 -435 -533 -59
rect -499 -435 -487 -59
rect -545 -447 -487 -435
rect -287 -59 -229 -47
rect -287 -435 -275 -59
rect -241 -435 -229 -59
rect -287 -447 -229 -435
rect -29 -59 29 -47
rect -29 -435 -17 -59
rect 17 -435 29 -59
rect -29 -447 29 -435
rect 229 -59 287 -47
rect 229 -435 241 -59
rect 275 -435 287 -59
rect 229 -447 287 -435
rect 487 -59 545 -47
rect 487 -435 499 -59
rect 533 -435 545 -59
rect 487 -447 545 -435
<< pdiffc >>
rect -533 130 -499 506
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect 499 130 533 506
rect -533 -435 -499 -59
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect 499 -435 533 -59
<< nsubdiff >>
rect -647 596 -551 630
rect 551 596 647 630
rect -647 -596 -613 596
rect 613 -596 647 596
rect -647 -630 647 -596
<< nsubdiffcont >>
rect -551 596 551 630
<< poly >>
rect -487 518 -287 544
rect -229 518 -29 544
rect 29 518 229 544
rect 287 518 487 544
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -47 -287 -21
rect -229 -47 -29 -21
rect 29 -47 229 -21
rect 287 -47 487 -21
rect -487 -494 -287 -447
rect -487 -528 -471 -494
rect -303 -528 -287 -494
rect -487 -544 -287 -528
rect -229 -494 -29 -447
rect -229 -528 -213 -494
rect -45 -528 -29 -494
rect -229 -544 -29 -528
rect 29 -494 229 -447
rect 29 -528 45 -494
rect 213 -528 229 -494
rect 29 -544 229 -528
rect 287 -494 487 -447
rect 287 -528 303 -494
rect 471 -528 487 -494
rect 287 -544 487 -528
<< polycont >>
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -528 -303 -494
rect -213 -528 -45 -494
rect 45 -528 213 -494
rect 303 -528 471 -494
<< locali >>
rect -647 -596 -613 630
rect -533 506 -499 522
rect -533 114 -499 130
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect 499 506 533 522
rect 499 114 533 130
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -533 -59 -499 -43
rect -533 -451 -499 -435
rect -275 -59 -241 -43
rect -275 -451 -241 -435
rect -17 -59 17 -43
rect -17 -451 17 -435
rect 241 -59 275 -43
rect 241 -451 275 -435
rect 499 -59 533 -43
rect 499 -451 533 -435
rect -487 -528 -471 -494
rect -303 -528 -287 -494
rect -229 -528 -213 -494
rect -45 -528 -29 -494
rect 29 -528 45 -494
rect 213 -528 229 -494
rect 287 -528 303 -494
rect 471 -528 487 -494
rect 613 -596 647 630
rect -647 -630 647 -596
<< viali >>
rect -613 596 -551 630
rect -551 596 551 630
rect 551 596 613 630
rect -533 130 -499 506
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect 499 130 533 506
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -533 -435 -499 -59
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect 499 -435 533 -59
rect -471 -528 -303 -494
rect -213 -528 -45 -494
rect 45 -528 213 -494
rect 303 -528 471 -494
<< metal1 >>
rect -625 630 625 636
rect -625 596 -613 630
rect 613 596 625 630
rect -625 590 625 596
rect -539 506 -493 518
rect -539 130 -533 506
rect -499 130 -493 506
rect -539 118 -493 130
rect -281 506 -235 518
rect -281 130 -275 506
rect -241 130 -235 506
rect -281 118 -235 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 235 506 281 518
rect 235 130 241 506
rect 275 130 281 506
rect 235 118 281 130
rect 493 506 539 518
rect 493 130 499 506
rect 533 130 539 506
rect 493 118 539 130
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect -539 -59 -493 -47
rect -539 -435 -533 -59
rect -499 -435 -493 -59
rect -539 -447 -493 -435
rect -281 -59 -235 -47
rect -281 -435 -275 -59
rect -241 -435 -235 -59
rect -281 -447 -235 -435
rect -23 -59 23 -47
rect -23 -435 -17 -59
rect 17 -435 23 -59
rect -23 -447 23 -435
rect 235 -59 281 -47
rect 235 -435 241 -59
rect 275 -435 281 -59
rect 235 -447 281 -435
rect 493 -59 539 -47
rect 493 -435 499 -59
rect 533 -435 539 -59
rect 493 -447 539 -435
rect -483 -494 -291 -488
rect -483 -528 -471 -494
rect -303 -528 -291 -494
rect -483 -534 -291 -528
rect -225 -494 -33 -488
rect -225 -528 -213 -494
rect -45 -528 -33 -494
rect -225 -534 -33 -528
rect 33 -494 225 -488
rect 33 -528 45 -494
rect 213 -528 225 -494
rect 33 -534 225 -528
rect 291 -494 483 -488
rect 291 -528 303 -494
rect 471 -528 483 -494
rect 291 -534 483 -528
<< properties >>
string FIXED_BBOX -630 -613 630 613
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
