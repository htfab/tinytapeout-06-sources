/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`define default_netname none

module tt_um_CDMA_Santiago (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
  //Instantiate cdma module
    cdma cdma_U1(  
        .clk_i(clk),
        .rst_i(~rst_n),
        .signal_i(ui_in[0]),
        .seed_i(ui_in[5:1]), 
        .receptor_i(ui_in[6]),
        .load_i(ui_in[7]),
        .cdma_o(uio_out[0]),
        .gold_o(uio_out[1]),
        .receptor_o(uio_out[2]),
        .led_o(uio_out[3])
    );
  // All output pins must be assigned. If not used, assign to 0.
    assign uio_oe = 8'b11111111;
    assign uo_out[7:0] = 8'b00000000;
    assign uio_out[7:4] = 4'b0000;
endmodule
