magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -683 -719 683 719
<< nmos >>
rect -487 109 -287 509
rect -229 109 -29 509
rect 29 109 229 509
rect 287 109 487 509
rect -487 -509 -287 -109
rect -229 -509 -29 -109
rect 29 -509 229 -109
rect 287 -509 487 -109
<< ndiff >>
rect -545 497 -487 509
rect -545 121 -533 497
rect -499 121 -487 497
rect -545 109 -487 121
rect -287 497 -229 509
rect -287 121 -275 497
rect -241 121 -229 497
rect -287 109 -229 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 229 497 287 509
rect 229 121 241 497
rect 275 121 287 497
rect 229 109 287 121
rect 487 497 545 509
rect 487 121 499 497
rect 533 121 545 497
rect 487 109 545 121
rect -545 -121 -487 -109
rect -545 -497 -533 -121
rect -499 -497 -487 -121
rect -545 -509 -487 -497
rect -287 -121 -229 -109
rect -287 -497 -275 -121
rect -241 -497 -229 -121
rect -287 -509 -229 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 229 -121 287 -109
rect 229 -497 241 -121
rect 275 -497 287 -121
rect 229 -509 287 -497
rect 487 -121 545 -109
rect 487 -497 499 -121
rect 533 -497 545 -121
rect 487 -509 545 -497
<< ndiffc >>
rect -533 121 -499 497
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect 499 121 533 497
rect -533 -497 -499 -121
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
rect 499 -497 533 -121
<< psubdiff >>
rect -647 649 -551 683
rect 551 649 647 683
rect -647 587 -613 649
rect 613 587 647 649
rect -647 -649 -613 -587
rect 613 -649 647 -587
rect -647 -683 647 -649
<< psubdiffcont >>
rect -551 649 551 683
rect -647 -587 -613 587
rect 613 -587 647 587
<< poly >>
rect -487 581 -287 597
rect -487 547 -471 581
rect -303 547 -287 581
rect -487 509 -287 547
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 509 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 509 229 547
rect 287 581 487 597
rect 287 547 303 581
rect 471 547 487 581
rect 287 509 487 547
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect -487 -547 -287 -509
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -487 -597 -287 -581
rect -229 -547 -29 -509
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -509
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
rect 287 -547 487 -509
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 287 -597 487 -581
<< polycont >>
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
<< locali >>
rect -647 587 -613 683
rect 613 587 647 683
rect -487 547 -471 581
rect -303 547 -287 581
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect 287 547 303 581
rect 471 547 487 581
rect -533 497 -499 513
rect -533 105 -499 121
rect -275 497 -241 513
rect -275 105 -241 121
rect -17 497 17 513
rect -17 105 17 121
rect 241 497 275 513
rect 241 105 275 121
rect 499 497 533 513
rect 499 105 533 121
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect -533 -121 -499 -105
rect -533 -513 -499 -497
rect -275 -121 -241 -105
rect -275 -513 -241 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 241 -121 275 -105
rect 241 -513 275 -497
rect 499 -121 533 -105
rect 499 -513 533 -497
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 287 -581 303 -547
rect 471 -581 487 -547
rect -647 -683 647 -649
<< viali >>
rect -613 649 -551 683
rect -551 649 551 683
rect 551 649 613 683
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect -533 330 -499 480
rect -275 138 -241 288
rect -17 330 17 480
rect 241 138 275 288
rect 499 330 533 480
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -647 -587 -613 -130
rect -533 -288 -499 -138
rect -275 -480 -241 -330
rect -17 -288 17 -138
rect 241 -480 275 -330
rect 499 -288 533 -138
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect -647 -649 -613 -587
rect 613 -587 647 -130
rect 613 -649 647 -587
<< metal1 >>
rect -625 683 625 689
rect -625 649 -613 683
rect 613 649 625 683
rect -625 643 625 649
rect -483 581 -291 587
rect -483 547 -471 581
rect -303 547 -291 581
rect -483 541 -291 547
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect 291 581 483 587
rect 291 547 303 581
rect 471 547 483 581
rect 291 541 483 547
rect -539 480 -493 492
rect -539 330 -533 480
rect -499 330 -493 480
rect -539 318 -493 330
rect -23 480 23 492
rect -23 330 -17 480
rect 17 330 23 480
rect -23 318 23 330
rect 493 480 539 492
rect 493 330 499 480
rect 533 330 539 480
rect 493 318 539 330
rect -281 288 -235 300
rect -281 138 -275 288
rect -241 138 -235 288
rect -281 126 -235 138
rect 235 288 281 300
rect 235 138 241 288
rect 275 138 281 288
rect 235 126 281 138
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect -653 -130 -607 -118
rect -653 -649 -647 -130
rect -613 -649 -607 -130
rect -539 -138 -493 -126
rect -539 -288 -533 -138
rect -499 -288 -493 -138
rect -539 -300 -493 -288
rect -23 -138 23 -126
rect -23 -288 -17 -138
rect 17 -288 23 -138
rect -23 -300 23 -288
rect 493 -138 539 -126
rect 493 -288 499 -138
rect 533 -288 539 -138
rect 493 -300 539 -288
rect 607 -130 653 -118
rect -281 -330 -235 -318
rect -281 -480 -275 -330
rect -241 -480 -235 -330
rect -281 -492 -235 -480
rect 235 -330 281 -318
rect 235 -480 241 -330
rect 275 -480 281 -330
rect 235 -492 281 -480
rect -483 -547 -291 -541
rect -483 -581 -471 -547
rect -303 -581 -291 -547
rect -483 -587 -291 -581
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
rect 291 -547 483 -541
rect 291 -581 303 -547
rect 471 -581 483 -547
rect 291 -587 483 -581
rect -653 -661 -607 -649
rect 607 -649 613 -130
rect 647 -649 653 -130
rect 607 -661 653 -649
<< properties >>
string FIXED_BBOX -630 -666 630 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
