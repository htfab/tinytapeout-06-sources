magic
tech sky130A
magscale 1 2
timestamp 1713334679
<< nwell >>
rect 690 -470 1610 -20
<< mvpsubdiff >>
rect 1446 -821 1470 -779
rect 1512 -821 1536 -779
<< mvnsubdiff >>
rect 1450 -128 1474 -86
rect 1516 -128 1540 -86
<< mvpsubdiffcont >>
rect 1470 -821 1512 -779
<< mvnsubdiffcont >>
rect 1474 -128 1516 -86
<< locali >>
rect 1458 -128 1474 -86
rect 1516 -128 1532 -86
rect 1454 -821 1470 -779
rect 1512 -821 1528 -779
<< viali >>
rect 1477 -125 1511 -91
rect 1475 -817 1509 -783
<< metal1 >>
rect 852 -55 1449 -17
rect 852 -70 890 -55
rect 690 -229 890 -70
rect 690 -267 968 -229
rect 690 -270 890 -267
rect 690 -475 890 -330
rect 1009 -450 1047 -89
rect 1167 -157 1205 -55
rect 1411 -85 1449 -55
rect 1167 -195 1248 -157
rect 1087 -375 1163 -337
rect 978 -475 1047 -450
rect 690 -513 1047 -475
rect 690 -530 890 -513
rect 978 -544 1047 -513
rect 690 -654 890 -590
rect 690 -692 968 -654
rect 690 -759 890 -692
rect 690 -790 891 -759
rect 1009 -774 1047 -544
rect 1125 -473 1163 -375
rect 1289 -441 1327 -89
rect 1411 -91 1523 -85
rect 1411 -125 1477 -91
rect 1511 -125 1523 -91
rect 1411 -127 1523 -125
rect 1465 -131 1523 -127
rect 1368 -330 1406 -251
rect 1368 -375 1640 -330
rect 1257 -473 1327 -441
rect 1125 -511 1327 -473
rect 1125 -595 1163 -511
rect 1257 -556 1327 -511
rect 1087 -633 1163 -595
rect 1173 -702 1252 -664
rect 853 -811 891 -790
rect 1173 -811 1211 -702
rect 1289 -774 1327 -556
rect 1405 -530 1640 -375
rect 1405 -595 1443 -530
rect 1367 -633 1443 -595
rect 1463 -781 1521 -777
rect 1410 -783 1521 -781
rect 1410 -811 1475 -783
rect 853 -817 1475 -811
rect 1509 -817 1521 -783
rect 853 -823 1521 -817
rect 853 -849 1450 -823
use sky130_fd_pr__nfet_g5v0d10v5_VNEAGC  sky130_fd_pr__nfet_g5v0d10v5_VNEAGC_0 cells
timestamp 1713334679
transform 1 0 1028 0 1 -652
box -108 -138 108 138
use sky130_fd_pr__nfet_g5v0d10v5_VNEAGC  sky130_fd_pr__nfet_g5v0d10v5_VNEAGC_2
timestamp 1713334679
transform 1 0 1308 0 1 -652
box -108 -138 108 138
use sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5  sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5_0 cells
timestamp 1713334679
transform 1 0 1308 0 1 -270
box -174 -200 174 200
use sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5  sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5_1
timestamp 1713334679
transform 1 0 1028 0 1 -270
box -174 -200 174 200
<< labels >>
flabel metal1 690 -790 890 -590 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 690 -530 890 -330 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 1440 -530 1640 -330 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 690 -270 890 -70 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
