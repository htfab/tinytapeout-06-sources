// This is the unpowered netlist.
module top (clk,
    rst_n,
    ui_in,
    uo_out);
 input clk;
 input rst_n;
 input [3:0] ui_in;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire \down_key.d ;
 wire \down_key.dff1 ;
 wire \down_key.dff2 ;
 wire \game.ballDirX ;
 wire \game.ballDirY ;
 wire \game.ballX[0] ;
 wire \game.ballX[1] ;
 wire \game.ballX[2] ;
 wire \game.ballX[3] ;
 wire \game.ballX[4] ;
 wire \game.ballX[5] ;
 wire \game.ballX[6] ;
 wire \game.ballX[7] ;
 wire \game.ballX[8] ;
 wire \game.ballY[0] ;
 wire \game.ballY[1] ;
 wire \game.ballY[2] ;
 wire \game.ballY[3] ;
 wire \game.ballY[4] ;
 wire \game.ballY[5] ;
 wire \game.ballY[6] ;
 wire \game.ballY[7] ;
 wire \game.blue ;
 wire \game.col0 ;
 wire \game.green ;
 wire \game.h[0] ;
 wire \game.h[1] ;
 wire \game.h[2] ;
 wire \game.h[3] ;
 wire \game.h[4] ;
 wire \game.h[5] ;
 wire \game.h[6] ;
 wire \game.h[7] ;
 wire \game.h[8] ;
 wire \game.h[9] ;
 wire \game.hit ;
 wire \game.hsync ;
 wire \game.inBallX ;
 wire \game.inBallY ;
 wire \game.inPaddle ;
 wire \game.new_game_n ;
 wire \game.offset[0] ;
 wire \game.offset[1] ;
 wire \game.offset[2] ;
 wire \game.offset[3] ;
 wire \game.offset[4] ;
 wire \game.paddle[0] ;
 wire \game.paddle[1] ;
 wire \game.paddle[2] ;
 wire \game.paddle[3] ;
 wire \game.paddle[4] ;
 wire \game.paddle[5] ;
 wire \game.paddle[6] ;
 wire \game.paddle[7] ;
 wire \game.paddle[8] ;
 wire \game.pause_n ;
 wire \game.red ;
 wire \game.row0 ;
 wire \game.speaker ;
 wire \game.up_key_n ;
 wire \game.v[0] ;
 wire \game.v[1] ;
 wire \game.v[2] ;
 wire \game.v[3] ;
 wire \game.v[4] ;
 wire \game.v[5] ;
 wire \game.v[6] ;
 wire \game.v[7] ;
 wire \game.v[8] ;
 wire \game.v[9] ;
 wire \game.vsync ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \new_game.d ;
 wire \new_game.dff1 ;
 wire \pause.d ;
 wire \pause.dff1 ;
 wire qb;
 wire qg;
 wire qr;
 wire \up_key.d ;
 wire \up_key.dff1 ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__or3_1 _0463_ (.A(\game.v[7] ),
    .B(\game.v[6] ),
    .C(\game.v[5] ),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _0464_ (.A(\game.v[4] ),
    .B(_0057_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_2 _0465_ (.A(\game.v[9] ),
    .X(_0059_));
 sky130_fd_sc_hd__or3_1 _0466_ (.A(\game.v[2] ),
    .B(\game.v[1] ),
    .C(\game.v[0] ),
    .X(_0060_));
 sky130_fd_sc_hd__or4_1 _0467_ (.A(_0059_),
    .B(\game.v[8] ),
    .C(\game.v[3] ),
    .D(_0060_),
    .X(_0061_));
 sky130_fd_sc_hd__nor2_1 _0468_ (.A(_0058_),
    .B(_0061_),
    .Y(\game.row0 ));
 sky130_fd_sc_hd__buf_2 _0469_ (.A(\game.h[0] ),
    .X(_0062_));
 sky130_fd_sc_hd__buf_2 _0470_ (.A(\game.h[5] ),
    .X(_0063_));
 sky130_fd_sc_hd__buf_2 _0471_ (.A(\game.h[1] ),
    .X(_0064_));
 sky130_fd_sc_hd__buf_2 _0472_ (.A(\game.h[2] ),
    .X(_0065_));
 sky130_fd_sc_hd__buf_2 _0473_ (.A(\game.h[4] ),
    .X(_0066_));
 sky130_fd_sc_hd__or4_1 _0474_ (.A(_0064_),
    .B(\game.h[3] ),
    .C(_0065_),
    .D(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__or2_1 _0475_ (.A(\game.h[7] ),
    .B(\game.h[8] ),
    .X(_0068_));
 sky130_fd_sc_hd__or3_1 _0476_ (.A(\game.h[6] ),
    .B(\game.h[9] ),
    .C(_0068_),
    .X(_0069_));
 sky130_fd_sc_hd__nor4_1 _0477_ (.A(_0062_),
    .B(_0063_),
    .C(_0067_),
    .D(_0069_),
    .Y(\game.col0 ));
 sky130_fd_sc_hd__or3b_1 _0478_ (.A(_0063_),
    .B(_0069_),
    .C_N(\game.inPaddle ),
    .X(_0070_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\game.v[1] ),
    .Y(_0071_));
 sky130_fd_sc_hd__or2_1 _0480_ (.A(\game.v[2] ),
    .B(\game.v[1] ),
    .X(_0072_));
 sky130_fd_sc_hd__nand2_1 _0481_ (.A(\game.v[3] ),
    .B(\game.v[2] ),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _0482_ (.A(\game.v[3] ),
    .Y(_0074_));
 sky130_fd_sc_hd__nor2_1 _0483_ (.A(\game.v[4] ),
    .B(_0074_),
    .Y(_0075_));
 sky130_fd_sc_hd__a221o_1 _0484_ (.A1(\game.v[4] ),
    .A2(_0071_),
    .B1(_0072_),
    .B2(_0073_),
    .C1(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__nand4_1 _0485_ (.A(_0064_),
    .B(\game.h[3] ),
    .C(_0065_),
    .D(_0066_),
    .Y(_0077_));
 sky130_fd_sc_hd__and3_1 _0486_ (.A(\game.v[8] ),
    .B(\game.v[7] ),
    .C(\game.v[6] ),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _0487_ (.A(_0063_),
    .B(\game.h[6] ),
    .X(_0079_));
 sky130_fd_sc_hd__o21ai_1 _0488_ (.A1(_0068_),
    .A2(_0079_),
    .B1(\game.h[9] ),
    .Y(_0080_));
 sky130_fd_sc_hd__or3_1 _0489_ (.A(\game.v[9] ),
    .B(\game.v[8] ),
    .C(_0057_),
    .X(_0081_));
 sky130_fd_sc_hd__and4bb_1 _0490_ (.A_N(_0059_),
    .B_N(_0078_),
    .C(_0080_),
    .D(_0081_),
    .X(_0082_));
 sky130_fd_sc_hd__a31o_1 _0491_ (.A1(_0067_),
    .A2(_0076_),
    .A3(_0077_),
    .B1(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_4 _0492_ (.A(\game.v[5] ),
    .X(_0084_));
 sky130_fd_sc_hd__a221o_1 _0493_ (.A1(\game.h[9] ),
    .A2(_0068_),
    .B1(_0078_),
    .B2(_0084_),
    .C1(_0059_),
    .X(_0085_));
 sky130_fd_sc_hd__a21oi_1 _0494_ (.A1(_0070_),
    .A2(_0083_),
    .B1(_0085_),
    .Y(\game.red ));
 sky130_fd_sc_hd__nand2_1 _0495_ (.A(\game.inBallY ),
    .B(net23),
    .Y(_0086_));
 sky130_fd_sc_hd__a21oi_1 _0496_ (.A1(_0082_),
    .A2(_0086_),
    .B1(_0085_),
    .Y(\game.green ));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(\game.v[2] ),
    .Y(_0087_));
 sky130_fd_sc_hd__and4b_1 _0498_ (.A_N(_0059_),
    .B(_0084_),
    .C(_0087_),
    .D(\game.v[1] ),
    .X(_0088_));
 sky130_fd_sc_hd__nand3_1 _0499_ (.A(_0078_),
    .B(_0075_),
    .C(_0088_),
    .Y(\game.vsync ));
 sky130_fd_sc_hd__or3_1 _0500_ (.A(_0063_),
    .B(_0066_),
    .C(\game.h[6] ),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_1 _0501_ (.A1(_0066_),
    .A2(_0079_),
    .B1(\game.h[8] ),
    .Y(_0090_));
 sky130_fd_sc_hd__nand4_1 _0502_ (.A(\game.h[7] ),
    .B(\game.h[9] ),
    .C(_0089_),
    .D(_0090_),
    .Y(\game.hsync ));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(net2),
    .Y(\pause.d ));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(net3),
    .Y(\new_game.d ));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(net4),
    .Y(\down_key.d ));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(net5),
    .Y(\up_key.d ));
 sky130_fd_sc_hd__or2_1 _0507_ (.A(\game.v[0] ),
    .B(_0062_),
    .X(_0091_));
 sky130_fd_sc_hd__nand2_1 _0508_ (.A(\game.v[0] ),
    .B(_0062_),
    .Y(_0092_));
 sky130_fd_sc_hd__or2b_1 _0509_ (.A(\game.offset[1] ),
    .B_N(\game.v[0] ),
    .X(_0093_));
 sky130_fd_sc_hd__or2b_1 _0510_ (.A(\game.v[0] ),
    .B_N(\game.offset[1] ),
    .X(_0094_));
 sky130_fd_sc_hd__or2b_1 _0511_ (.A(\game.h[3] ),
    .B_N(\game.offset[4] ),
    .X(_0095_));
 sky130_fd_sc_hd__or2b_1 _0512_ (.A(\game.h[1] ),
    .B_N(\game.offset[2] ),
    .X(_0096_));
 sky130_fd_sc_hd__or2b_1 _0513_ (.A(_0062_),
    .B_N(\game.offset[1] ),
    .X(_0097_));
 sky130_fd_sc_hd__and2b_1 _0514_ (.A_N(\game.offset[2] ),
    .B(_0064_),
    .X(_0098_));
 sky130_fd_sc_hd__a21oi_1 _0515_ (.A1(_0096_),
    .A2(_0097_),
    .B1(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__and2b_1 _0516_ (.A_N(_0065_),
    .B(\game.offset[3] ),
    .X(_0100_));
 sky130_fd_sc_hd__or2b_1 _0517_ (.A(\game.offset[3] ),
    .B_N(_0065_),
    .X(_0101_));
 sky130_fd_sc_hd__o21ai_1 _0518_ (.A1(_0099_),
    .A2(_0100_),
    .B1(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__and2b_1 _0519_ (.A_N(\game.offset[4] ),
    .B(\game.h[3] ),
    .X(_0103_));
 sky130_fd_sc_hd__a21oi_1 _0520_ (.A1(_0095_),
    .A2(_0102_),
    .B1(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__xnor2_1 _0521_ (.A(_0066_),
    .B(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_1 _0522_ (.A(_0074_),
    .B(\game.offset[4] ),
    .Y(_0106_));
 sky130_fd_sc_hd__or2b_1 _0523_ (.A(\game.v[1] ),
    .B_N(\game.offset[2] ),
    .X(_0107_));
 sky130_fd_sc_hd__and2b_1 _0524_ (.A_N(\game.offset[2] ),
    .B(\game.v[1] ),
    .X(_0108_));
 sky130_fd_sc_hd__a21o_1 _0525_ (.A1(_0107_),
    .A2(_0094_),
    .B1(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_1 _0526_ (.A(_0087_),
    .B(\game.offset[3] ),
    .Y(_0110_));
 sky130_fd_sc_hd__nor2_1 _0527_ (.A(_0087_),
    .B(\game.offset[3] ),
    .Y(_0111_));
 sky130_fd_sc_hd__a21o_1 _0528_ (.A1(_0109_),
    .A2(_0110_),
    .B1(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__nor2_1 _0529_ (.A(_0074_),
    .B(\game.offset[4] ),
    .Y(_0113_));
 sky130_fd_sc_hd__a21oi_1 _0530_ (.A1(_0106_),
    .A2(_0112_),
    .B1(_0113_),
    .Y(_0114_));
 sky130_fd_sc_hd__xnor2_1 _0531_ (.A(\game.v[4] ),
    .B(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__xnor2_1 _0532_ (.A(_0105_),
    .B(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__a221oi_1 _0533_ (.A1(_0091_),
    .A2(_0092_),
    .B1(_0093_),
    .B2(_0094_),
    .C1(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__xor2_1 _0534_ (.A(\game.v[2] ),
    .B(_0065_),
    .X(_0118_));
 sky130_fd_sc_hd__xnor2_1 _0535_ (.A(_0099_),
    .B(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__xnor2_1 _0536_ (.A(_0109_),
    .B(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__and2b_1 _0537_ (.A_N(_0103_),
    .B(_0095_),
    .X(_0121_));
 sky130_fd_sc_hd__xnor2_1 _0538_ (.A(_0102_),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__and2b_1 _0539_ (.A_N(_0113_),
    .B(_0106_),
    .X(_0123_));
 sky130_fd_sc_hd__xnor2_1 _0540_ (.A(_0112_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__xor2_1 _0541_ (.A(_0122_),
    .B(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__xnor2_1 _0542_ (.A(_0120_),
    .B(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__and4_1 _0543_ (.A(_0116_),
    .B(_0091_),
    .C(_0092_),
    .D(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__or2b_1 _0544_ (.A(_0116_),
    .B_N(_0126_),
    .X(_0128_));
 sky130_fd_sc_hd__o211a_1 _0545_ (.A1(_0085_),
    .A2(_0070_),
    .B1(_0082_),
    .C1(_0086_),
    .X(_0129_));
 sky130_fd_sc_hd__o211a_1 _0546_ (.A1(_0117_),
    .A2(_0127_),
    .B1(_0128_),
    .C1(_0129_),
    .X(\game.blue ));
 sky130_fd_sc_hd__or2_1 _0547_ (.A(\game.ballX[3] ),
    .B(\game.ballX[4] ),
    .X(_0130_));
 sky130_fd_sc_hd__nor2_1 _0548_ (.A(\game.ballX[6] ),
    .B(\game.ballX[7] ),
    .Y(_0131_));
 sky130_fd_sc_hd__a21bo_1 _0549_ (.A1(\game.ballX[5] ),
    .A2(_0130_),
    .B1_N(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__and2_1 _0550_ (.A(\game.ballY[3] ),
    .B(\game.ballY[4] ),
    .X(_0133_));
 sky130_fd_sc_hd__o211a_1 _0551_ (.A1(\game.ballY[5] ),
    .A2(_0133_),
    .B1(\game.ballY[7] ),
    .C1(\game.ballY[6] ),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _0552_ (.A(\game.ballY[4] ),
    .B(\game.ballY[5] ),
    .X(_0135_));
 sky130_fd_sc_hd__nor3_1 _0553_ (.A(\game.ballY[6] ),
    .B(\game.ballY[7] ),
    .C(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__a211o_1 _0554_ (.A1(\game.ballX[8] ),
    .A2(_0132_),
    .B1(_0134_),
    .C1(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _0555_ (.A1(_0084_),
    .A2(\game.hit ),
    .B1(_0137_),
    .B2(\game.v[6] ),
    .X(\game.speaker ));
 sky130_fd_sc_hd__buf_2 _0556_ (.A(net1),
    .X(_0138_));
 sky130_fd_sc_hd__nor2_1 _0557_ (.A(\game.h[5] ),
    .B(\game.h[6] ),
    .Y(_0139_));
 sky130_fd_sc_hd__and4_2 _0558_ (.A(\game.h[1] ),
    .B(\game.h[0] ),
    .C(\game.h[3] ),
    .D(\game.h[2] ),
    .X(_0140_));
 sky130_fd_sc_hd__and3b_1 _0559_ (.A_N(\game.h[7] ),
    .B(\game.h[9] ),
    .C(\game.h[8] ),
    .X(_0141_));
 sky130_fd_sc_hd__and4_2 _0560_ (.A(\game.h[4] ),
    .B(_0139_),
    .C(_0140_),
    .D(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__or4b_1 _0561_ (.A(\game.v[8] ),
    .B(\game.v[1] ),
    .C(\game.v[0] ),
    .D_N(\game.v[9] ),
    .X(_0143_));
 sky130_fd_sc_hd__nor3_1 _0562_ (.A(_0058_),
    .B(_0073_),
    .C(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__and3_2 _0563_ (.A(\game.pause_n ),
    .B(_0142_),
    .C(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__or2_1 _0564_ (.A(\game.offset[0] ),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_4 _0565_ (.A(_0145_),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_1 _0566_ (.A(\game.offset[0] ),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__and3_1 _0567_ (.A(_0138_),
    .B(_0146_),
    .C(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _0568_ (.A(_0149_),
    .X(_0000_));
 sky130_fd_sc_hd__and3_1 _0569_ (.A(\game.offset[1] ),
    .B(\game.offset[0] ),
    .C(_0145_),
    .X(_0150_));
 sky130_fd_sc_hd__nand4_2 _0570_ (.A(\game.h[4] ),
    .B(_0139_),
    .C(_0140_),
    .D(_0141_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor4_1 _0571_ (.A(_0058_),
    .B(_0073_),
    .C(_0151_),
    .D(_0143_),
    .Y(_0152_));
 sky130_fd_sc_hd__a31o_1 _0572_ (.A1(\game.offset[0] ),
    .A2(\game.pause_n ),
    .A3(_0152_),
    .B1(\game.offset[1] ),
    .X(_0153_));
 sky130_fd_sc_hd__and3b_1 _0573_ (.A_N(_0150_),
    .B(_0138_),
    .C(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _0574_ (.A(_0154_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _0575_ (.A(\game.offset[2] ),
    .B(_0150_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _0576_ (.A(\game.offset[2] ),
    .B(_0150_),
    .Y(_0156_));
 sky130_fd_sc_hd__and3_1 _0577_ (.A(_0138_),
    .B(_0155_),
    .C(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _0578_ (.A(_0157_),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _0579_ (.A(\game.offset[3] ),
    .B(\game.offset[2] ),
    .C(_0150_),
    .X(_0158_));
 sky130_fd_sc_hd__a21o_1 _0580_ (.A1(\game.offset[2] ),
    .A2(_0150_),
    .B1(\game.offset[3] ),
    .X(_0159_));
 sky130_fd_sc_hd__and3b_1 _0581_ (.A_N(_0158_),
    .B(_0138_),
    .C(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0582_ (.A(_0160_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_4 _0583_ (.A(net1),
    .X(_0161_));
 sky130_fd_sc_hd__o21ai_1 _0584_ (.A1(net12),
    .A2(_0158_),
    .B1(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__a21oi_1 _0585_ (.A1(net12),
    .A2(_0158_),
    .B1(_0162_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_2 _0586_ (.A(\game.pause_n ),
    .B(net6),
    .Y(_0163_));
 sky130_fd_sc_hd__a21oi_1 _0587_ (.A1(\game.paddle[7] ),
    .A2(\game.paddle[8] ),
    .B1(\down_key.dff2 ),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _0588_ (.A(\game.up_key_n ),
    .Y(_0165_));
 sky130_fd_sc_hd__o41a_1 _0589_ (.A1(\game.paddle[7] ),
    .A2(\game.paddle[6] ),
    .A3(\game.paddle[5] ),
    .A4(\game.paddle[8] ),
    .B1(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_1 _0590_ (.A(_0164_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__nor2_2 _0591_ (.A(_0163_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__or2_1 _0592_ (.A(\game.new_game_n ),
    .B(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__and3_1 _0593_ (.A(net19),
    .B(_0138_),
    .C(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0594_ (.A(_0170_),
    .X(_0005_));
 sky130_fd_sc_hd__o21a_1 _0595_ (.A1(_0163_),
    .A2(_0167_),
    .B1(\game.new_game_n ),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(_0168_),
    .A1(_0171_),
    .S(\game.paddle[1] ),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _0597_ (.A(_0161_),
    .B(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _0598_ (.A(_0173_),
    .X(_0006_));
 sky130_fd_sc_hd__a21o_2 _0599_ (.A1(\game.paddle[7] ),
    .A2(\game.paddle[8] ),
    .B1(\down_key.dff2 ),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _0600_ (.A(_0174_),
    .B(_0166_),
    .X(_0175_));
 sky130_fd_sc_hd__xor2_1 _0601_ (.A(\game.paddle[2] ),
    .B(\game.paddle[1] ),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(_0164_),
    .A1(_0175_),
    .S(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__o2bb2a_1 _0603_ (.A1_N(_0145_),
    .A2_N(_0177_),
    .B1(_0168_),
    .B2(\game.paddle[2] ),
    .X(_0178_));
 sky130_fd_sc_hd__and3_1 _0604_ (.A(_0138_),
    .B(_0169_),
    .C(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0605_ (.A(_0179_),
    .X(_0007_));
 sky130_fd_sc_hd__o21ai_1 _0606_ (.A1(\game.paddle[2] ),
    .A2(\game.paddle[1] ),
    .B1(\game.paddle[3] ),
    .Y(_0180_));
 sky130_fd_sc_hd__or3_2 _0607_ (.A(\game.paddle[3] ),
    .B(\game.paddle[2] ),
    .C(\game.paddle[1] ),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _0608_ (.A(_0180_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__a31oi_2 _0609_ (.A1(\game.paddle[3] ),
    .A2(\game.paddle[2] ),
    .A3(\game.paddle[1] ),
    .B1(_0174_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21o_1 _0610_ (.A1(\game.paddle[2] ),
    .A2(\game.paddle[1] ),
    .B1(\game.paddle[3] ),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _0611_ (.A1(_0175_),
    .A2(_0182_),
    .B1(_0183_),
    .B2(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _0612_ (.A1(\game.paddle[3] ),
    .A2(_0171_),
    .B1(_0185_),
    .B2(_0147_),
    .X(_0186_));
 sky130_fd_sc_hd__and2_1 _0613_ (.A(_0161_),
    .B(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _0614_ (.A(_0187_),
    .X(_0008_));
 sky130_fd_sc_hd__a211o_1 _0615_ (.A1(_0174_),
    .A2(_0181_),
    .B1(_0183_),
    .C1(\game.paddle[4] ),
    .X(_0188_));
 sky130_fd_sc_hd__a31o_1 _0616_ (.A1(_0174_),
    .A2(_0166_),
    .A3(_0181_),
    .B1(_0183_),
    .X(_0189_));
 sky130_fd_sc_hd__a2bb2o_1 _0617_ (.A1_N(_0167_),
    .A2_N(_0188_),
    .B1(_0189_),
    .B2(\game.paddle[4] ),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_1 _0618_ (.A1(\game.paddle[4] ),
    .A2(_0171_),
    .B1(_0190_),
    .B2(_0147_),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _0619_ (.A(_0161_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0620_ (.A(_0192_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _0621_ (.A(net1),
    .X(_0193_));
 sky130_fd_sc_hd__and4_1 _0622_ (.A(\game.paddle[4] ),
    .B(\game.paddle[3] ),
    .C(\game.paddle[2] ),
    .D(\game.paddle[1] ),
    .X(_0194_));
 sky130_fd_sc_hd__and2_1 _0623_ (.A(\game.paddle[5] ),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _0624_ (.A(_0174_),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__nor2_1 _0625_ (.A(\game.paddle[5] ),
    .B(_0194_),
    .Y(_0197_));
 sky130_fd_sc_hd__or3_1 _0626_ (.A(\game.paddle[4] ),
    .B(\game.paddle[5] ),
    .C(_0181_),
    .X(_0198_));
 sky130_fd_sc_hd__o21ai_1 _0627_ (.A1(\game.paddle[4] ),
    .A2(_0181_),
    .B1(\game.paddle[5] ),
    .Y(_0199_));
 sky130_fd_sc_hd__a21bo_1 _0628_ (.A1(_0198_),
    .A2(_0199_),
    .B1_N(_0175_),
    .X(_0200_));
 sky130_fd_sc_hd__o21ai_1 _0629_ (.A1(_0196_),
    .A2(_0197_),
    .B1(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__a22o_1 _0630_ (.A1(\game.paddle[5] ),
    .A2(_0171_),
    .B1(_0201_),
    .B2(_0147_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _0631_ (.A(_0193_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(_0203_),
    .X(_0010_));
 sky130_fd_sc_hd__inv_2 _0633_ (.A(net17),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _0634_ (.A(_0174_),
    .B(_0198_),
    .Y(_0205_));
 sky130_fd_sc_hd__and3_1 _0635_ (.A(_0168_),
    .B(_0196_),
    .C(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__a21oi_1 _0636_ (.A1(_0204_),
    .A2(_0169_),
    .B1(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(net1),
    .Y(_0208_));
 sky130_fd_sc_hd__clkbuf_4 _0638_ (.A(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__a211o_1 _0639_ (.A1(_0204_),
    .A2(_0206_),
    .B1(_0207_),
    .C1(_0209_),
    .X(_0011_));
 sky130_fd_sc_hd__o21ai_1 _0640_ (.A1(\game.new_game_n ),
    .A2(_0168_),
    .B1(\game.paddle[7] ),
    .Y(_0210_));
 sky130_fd_sc_hd__or2_1 _0641_ (.A(\game.paddle[6] ),
    .B(_0198_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_4 _0642_ (.A(_0163_),
    .X(_0212_));
 sky130_fd_sc_hd__a21oi_1 _0643_ (.A1(\game.paddle[6] ),
    .A2(_0195_),
    .B1(_0174_),
    .Y(_0213_));
 sky130_fd_sc_hd__a2111o_1 _0644_ (.A1(_0174_),
    .A2(_0211_),
    .B1(_0167_),
    .C1(_0212_),
    .D1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0645_ (.A0(\game.paddle[7] ),
    .A1(_0210_),
    .S(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nor2_1 _0646_ (.A(_0209_),
    .B(_0215_),
    .Y(_0012_));
 sky130_fd_sc_hd__a31o_1 _0647_ (.A1(\game.paddle[7] ),
    .A2(\game.paddle[6] ),
    .A3(_0195_),
    .B1(_0174_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ai_1 _0648_ (.A1(\game.paddle[7] ),
    .A2(_0211_),
    .B1(_0174_),
    .Y(_0217_));
 sky130_fd_sc_hd__a41o_1 _0649_ (.A1(\game.paddle[8] ),
    .A2(_0168_),
    .A3(_0216_),
    .A4(_0217_),
    .B1(_0208_),
    .X(_0218_));
 sky130_fd_sc_hd__a32o_1 _0650_ (.A1(_0168_),
    .A2(_0216_),
    .A3(_0217_),
    .B1(_0169_),
    .B2(\game.paddle[8] ),
    .X(_0219_));
 sky130_fd_sc_hd__and2b_1 _0651_ (.A_N(_0218_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _0652_ (.A(_0220_),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _0653_ (.A(\game.ballY[0] ),
    .Y(_0221_));
 sky130_fd_sc_hd__and2_2 _0654_ (.A(\game.new_game_n ),
    .B(_0163_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_4 _0655_ (.A(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _0656_ (.A(_0221_),
    .B(_0212_),
    .Y(_0224_));
 sky130_fd_sc_hd__o211a_1 _0657_ (.A1(_0221_),
    .A2(_0223_),
    .B1(_0224_),
    .C1(_0161_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _0658_ (.A(\game.ballDirY ),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_2 _0659_ (.A(_0225_),
    .B(\game.ballY[1] ),
    .Y(_0226_));
 sky130_fd_sc_hd__xnor2_1 _0660_ (.A(\game.ballY[0] ),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__a22o_1 _0661_ (.A1(\game.ballY[1] ),
    .A2(_0223_),
    .B1(_0227_),
    .B2(_0147_),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _0662_ (.A(_0193_),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _0663_ (.A(_0229_),
    .X(_0015_));
 sky130_fd_sc_hd__nand2_1 _0664_ (.A(_0225_),
    .B(\game.ballY[1] ),
    .Y(_0230_));
 sky130_fd_sc_hd__o21ai_2 _0665_ (.A1(_0221_),
    .A2(_0226_),
    .B1(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__and2b_1 _0666_ (.A_N(\game.ballY[2] ),
    .B(_0225_),
    .X(_0232_));
 sky130_fd_sc_hd__and2b_1 _0667_ (.A_N(_0225_),
    .B(\game.ballY[2] ),
    .X(_0233_));
 sky130_fd_sc_hd__nor2_1 _0668_ (.A(_0232_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__xor2_1 _0669_ (.A(_0231_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _0670_ (.A1(\game.ballY[2] ),
    .A2(_0223_),
    .B1(_0235_),
    .B2(_0147_),
    .X(_0236_));
 sky130_fd_sc_hd__and2_1 _0671_ (.A(_0193_),
    .B(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0237_),
    .X(_0016_));
 sky130_fd_sc_hd__xor2_1 _0673_ (.A(_0225_),
    .B(\game.ballY[3] ),
    .X(_0238_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__a21oi_1 _0675_ (.A1(_0231_),
    .A2(_0234_),
    .B1(_0233_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_1 _0676_ (.A(_0239_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__a22o_1 _0677_ (.A1(\game.ballY[3] ),
    .A2(_0223_),
    .B1(_0241_),
    .B2(_0147_),
    .X(_0242_));
 sky130_fd_sc_hd__and2_1 _0678_ (.A(_0193_),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_1 _0679_ (.A(_0243_),
    .X(_0017_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(_0225_),
    .Y(_0244_));
 sky130_fd_sc_hd__o21a_1 _0681_ (.A1(\game.ballY[2] ),
    .A2(\game.ballY[3] ),
    .B1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__a31o_1 _0682_ (.A1(_0231_),
    .A2(_0234_),
    .A3(_0239_),
    .B1(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_1 _0683_ (.A(_0244_),
    .B(\game.ballY[4] ),
    .Y(_0247_));
 sky130_fd_sc_hd__and2_1 _0684_ (.A(_0244_),
    .B(\game.ballY[4] ),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _0685_ (.A(_0247_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__xor2_1 _0686_ (.A(_0246_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _0687_ (.A1(\game.ballY[4] ),
    .A2(_0223_),
    .B1(_0250_),
    .B2(_0147_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_1 _0688_ (.A(_0193_),
    .B(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _0689_ (.A(_0252_),
    .X(_0018_));
 sky130_fd_sc_hd__a21oi_1 _0690_ (.A1(_0246_),
    .A2(_0249_),
    .B1(_0248_),
    .Y(_0253_));
 sky130_fd_sc_hd__xnor2_1 _0691_ (.A(_0225_),
    .B(\game.ballY[5] ),
    .Y(_0254_));
 sky130_fd_sc_hd__a21oi_1 _0692_ (.A1(_0253_),
    .A2(_0254_),
    .B1(_0212_),
    .Y(_0255_));
 sky130_fd_sc_hd__or2_1 _0693_ (.A(_0253_),
    .B(_0254_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _0694_ (.A(\game.new_game_n ),
    .B(_0212_),
    .Y(_0257_));
 sky130_fd_sc_hd__o2bb2a_1 _0695_ (.A1_N(_0255_),
    .A2_N(_0256_),
    .B1(_0257_),
    .B2(\game.ballY[5] ),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _0696_ (.A(_0209_),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0259_),
    .X(_0019_));
 sky130_fd_sc_hd__and3_1 _0698_ (.A(\game.new_game_n ),
    .B(\game.ballY[6] ),
    .C(_0212_),
    .X(_0260_));
 sky130_fd_sc_hd__xnor2_1 _0699_ (.A(_0225_),
    .B(\game.ballY[6] ),
    .Y(_0261_));
 sky130_fd_sc_hd__a32o_1 _0700_ (.A1(_0246_),
    .A2(_0249_),
    .A3(_0254_),
    .B1(_0135_),
    .B2(_0244_),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _0701_ (.A(_0261_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(_0261_),
    .B(_0262_),
    .Y(_0264_));
 sky130_fd_sc_hd__and3_1 _0703_ (.A(_0147_),
    .B(_0263_),
    .C(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__o21a_1 _0704_ (.A1(_0260_),
    .A2(_0265_),
    .B1(_0161_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _0705_ (.A(net13),
    .B(_0223_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _0706_ (.A(_0244_),
    .B(\game.ballY[6] ),
    .Y(_0267_));
 sky130_fd_sc_hd__or2_1 _0707_ (.A(_0225_),
    .B(\game.ballY[7] ),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_1 _0708_ (.A(_0225_),
    .B(\game.ballY[7] ),
    .Y(_0269_));
 sky130_fd_sc_hd__and4_1 _0709_ (.A(_0267_),
    .B(_0264_),
    .C(_0268_),
    .D(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _0710_ (.A1(_0267_),
    .A2(_0264_),
    .B1(_0268_),
    .B2(_0269_),
    .X(_0271_));
 sky130_fd_sc_hd__or3b_1 _0711_ (.A(_0270_),
    .B(_0212_),
    .C_N(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__a21oi_1 _0712_ (.A1(_0266_),
    .A2(_0272_),
    .B1(_0209_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(\game.ballX[0] ),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _0714_ (.A(_0273_),
    .B(_0212_),
    .Y(_0274_));
 sky130_fd_sc_hd__o211a_1 _0715_ (.A1(_0273_),
    .A2(_0223_),
    .B1(_0274_),
    .C1(_0161_),
    .X(_0022_));
 sky130_fd_sc_hd__xnor2_1 _0716_ (.A(\game.ballDirX ),
    .B(\game.ballX[1] ),
    .Y(_0275_));
 sky130_fd_sc_hd__xnor2_1 _0717_ (.A(\game.ballX[0] ),
    .B(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__a22o_1 _0718_ (.A1(\game.ballX[1] ),
    .A2(_0222_),
    .B1(_0276_),
    .B2(_0147_),
    .X(_0277_));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(_0193_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_1 _0720_ (.A(_0278_),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _0721_ (.A(\game.ballDirX ),
    .B(\game.ballX[1] ),
    .Y(_0279_));
 sky130_fd_sc_hd__o21ai_2 _0722_ (.A1(_0273_),
    .A2(_0275_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__and2b_1 _0723_ (.A_N(\game.ballX[2] ),
    .B(\game.ballDirX ),
    .X(_0281_));
 sky130_fd_sc_hd__and2b_1 _0724_ (.A_N(\game.ballDirX ),
    .B(\game.ballX[2] ),
    .X(_0282_));
 sky130_fd_sc_hd__nor2_1 _0725_ (.A(_0281_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__xor2_1 _0726_ (.A(_0280_),
    .B(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(\game.ballX[2] ),
    .A2(_0222_),
    .B1(_0284_),
    .B2(_0145_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_1 _0728_ (.A(_0193_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _0729_ (.A(_0286_),
    .X(_0024_));
 sky130_fd_sc_hd__xnor2_1 _0730_ (.A(\game.ballDirX ),
    .B(\game.ballX[3] ),
    .Y(_0287_));
 sky130_fd_sc_hd__a21oi_1 _0731_ (.A1(_0280_),
    .A2(_0283_),
    .B1(_0282_),
    .Y(_0288_));
 sky130_fd_sc_hd__xnor2_1 _0732_ (.A(_0287_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(\game.ballX[3] ),
    .A2(_0222_),
    .B1(_0289_),
    .B2(_0145_),
    .X(_0290_));
 sky130_fd_sc_hd__and2_1 _0734_ (.A(_0193_),
    .B(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0291_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_2 _0736_ (.A(\game.ballX[4] ),
    .X(_0292_));
 sky130_fd_sc_hd__o21ba_1 _0737_ (.A1(\game.ballX[2] ),
    .A2(\game.ballX[3] ),
    .B1_N(\game.ballDirX ),
    .X(_0293_));
 sky130_fd_sc_hd__a31o_1 _0738_ (.A1(_0280_),
    .A2(_0283_),
    .A3(_0287_),
    .B1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_4 _0739_ (.A(\game.ballDirX ),
    .X(_0295_));
 sky130_fd_sc_hd__and2b_1 _0740_ (.A_N(_0292_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__and2b_1 _0741_ (.A_N(_0295_),
    .B(_0292_),
    .X(_0297_));
 sky130_fd_sc_hd__nor2_1 _0742_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__xor2_1 _0743_ (.A(_0294_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__a22o_1 _0744_ (.A1(_0292_),
    .A2(_0222_),
    .B1(_0299_),
    .B2(_0145_),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _0745_ (.A(_0193_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0746_ (.A(_0301_),
    .X(_0026_));
 sky130_fd_sc_hd__xor2_1 _0747_ (.A(_0295_),
    .B(\game.ballX[5] ),
    .X(_0302_));
 sky130_fd_sc_hd__a21o_1 _0748_ (.A1(_0294_),
    .A2(_0298_),
    .B1(_0297_),
    .X(_0303_));
 sky130_fd_sc_hd__nor2_1 _0749_ (.A(_0302_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__a21o_1 _0750_ (.A1(_0302_),
    .A2(_0303_),
    .B1(_0212_),
    .X(_0305_));
 sky130_fd_sc_hd__o22a_1 _0751_ (.A1(\game.ballX[5] ),
    .A2(_0257_),
    .B1(_0304_),
    .B2(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _0752_ (.A(_0209_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0307_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(net14),
    .B(_0223_),
    .Y(_0308_));
 sky130_fd_sc_hd__or2b_1 _0755_ (.A(\game.ballX[6] ),
    .B_N(_0295_),
    .X(_0309_));
 sky130_fd_sc_hd__or2b_1 _0756_ (.A(_0295_),
    .B_N(\game.ballX[6] ),
    .X(_0310_));
 sky130_fd_sc_hd__nand2_1 _0757_ (.A(_0309_),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__or4b_1 _0758_ (.A(_0296_),
    .B(_0302_),
    .C(_0297_),
    .D_N(_0294_),
    .X(_0312_));
 sky130_fd_sc_hd__o21bai_1 _0759_ (.A1(_0292_),
    .A2(\game.ballX[5] ),
    .B1_N(_0295_),
    .Y(_0313_));
 sky130_fd_sc_hd__and3_1 _0760_ (.A(_0311_),
    .B(_0312_),
    .C(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__a21o_1 _0761_ (.A1(_0312_),
    .A2(_0313_),
    .B1(_0311_),
    .X(_0315_));
 sky130_fd_sc_hd__or3b_1 _0762_ (.A(_0212_),
    .B(_0314_),
    .C_N(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__a21oi_1 _0763_ (.A1(_0308_),
    .A2(_0316_),
    .B1(_0209_),
    .Y(_0028_));
 sky130_fd_sc_hd__xor2_1 _0764_ (.A(_0295_),
    .B(\game.ballX[7] ),
    .X(_0317_));
 sky130_fd_sc_hd__a21oi_1 _0765_ (.A1(_0310_),
    .A2(_0315_),
    .B1(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__a31o_1 _0766_ (.A1(_0310_),
    .A2(_0315_),
    .A3(_0317_),
    .B1(_0212_),
    .X(_0319_));
 sky130_fd_sc_hd__o2bb2a_1 _0767_ (.A1_N(\game.ballX[7] ),
    .A2_N(_0223_),
    .B1(_0318_),
    .B2(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__nor2_1 _0768_ (.A(_0209_),
    .B(_0320_),
    .Y(_0029_));
 sky130_fd_sc_hd__or3_1 _0769_ (.A(_0311_),
    .B(_0312_),
    .C(_0317_),
    .X(_0321_));
 sky130_fd_sc_hd__o21a_1 _0770_ (.A1(_0295_),
    .A2(_0131_),
    .B1(_0313_),
    .X(_0322_));
 sky130_fd_sc_hd__xor2_1 _0771_ (.A(_0295_),
    .B(\game.ballX[8] ),
    .X(_0323_));
 sky130_fd_sc_hd__a21oi_1 _0772_ (.A1(_0321_),
    .A2(_0322_),
    .B1(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a31o_1 _0773_ (.A1(_0321_),
    .A2(_0322_),
    .A3(_0323_),
    .B1(_0163_),
    .X(_0325_));
 sky130_fd_sc_hd__a2bb2o_1 _0774_ (.A1_N(_0324_),
    .A2_N(_0325_),
    .B1(\game.ballX[8] ),
    .B2(_0223_),
    .X(_0326_));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(_0193_),
    .B(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0776_ (.A(_0327_),
    .X(_0030_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(_0084_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_1 _0778_ (.A(\game.v[0] ),
    .B(\game.paddle[0] ),
    .X(_0329_));
 sky130_fd_sc_hd__a221o_1 _0779_ (.A1(_0328_),
    .A2(\game.paddle[5] ),
    .B1(\game.paddle[2] ),
    .B2(_0087_),
    .C1(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(\game.paddle[3] ),
    .Y(_0331_));
 sky130_fd_sc_hd__o22a_1 _0781_ (.A1(_0328_),
    .A2(\game.paddle[5] ),
    .B1(\game.paddle[2] ),
    .B2(_0087_),
    .X(_0332_));
 sky130_fd_sc_hd__o221ai_1 _0782_ (.A1(\game.v[3] ),
    .A2(_0331_),
    .B1(\game.paddle[1] ),
    .B2(_0071_),
    .C1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__xor2_1 _0783_ (.A(\game.v[4] ),
    .B(\game.paddle[4] ),
    .X(_0334_));
 sky130_fd_sc_hd__a221o_1 _0784_ (.A1(\game.v[3] ),
    .A2(_0331_),
    .B1(\game.paddle[1] ),
    .B2(_0071_),
    .C1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__or4_1 _0785_ (.A(_0151_),
    .B(_0330_),
    .C(_0333_),
    .D(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__or2b_1 _0786_ (.A(\game.paddle[6] ),
    .B_N(\game.v[6] ),
    .X(_0337_));
 sky130_fd_sc_hd__or2b_1 _0787_ (.A(\game.v[6] ),
    .B_N(\game.paddle[6] ),
    .X(_0338_));
 sky130_fd_sc_hd__xor2_1 _0788_ (.A(\game.v[7] ),
    .B(\game.paddle[7] ),
    .X(_0339_));
 sky130_fd_sc_hd__xor2_1 _0789_ (.A(\game.v[8] ),
    .B(\game.paddle[8] ),
    .X(_0340_));
 sky130_fd_sc_hd__nor2_1 _0790_ (.A(_0339_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__and4b_1 _0791_ (.A_N(_0336_),
    .B(_0337_),
    .C(_0338_),
    .D(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _0792_ (.A(_0070_),
    .B(_0086_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21o_1 _0793_ (.A1(\game.new_game_n ),
    .A2(\game.hit ),
    .B1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__and3b_1 _0794_ (.A_N(_0342_),
    .B(_0344_),
    .C(net1),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0795_ (.A(_0345_),
    .X(_0031_));
 sky130_fd_sc_hd__and4_1 _0796_ (.A(\game.ballX[3] ),
    .B(_0292_),
    .C(\game.ballX[5] ),
    .D(\game.ballX[6] ),
    .X(_0346_));
 sky130_fd_sc_hd__xnor2_1 _0797_ (.A(\game.h[8] ),
    .B(\game.ballX[7] ),
    .Y(_0347_));
 sky130_fd_sc_hd__xnor2_1 _0798_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_1 _0799_ (.A(\game.h[9] ),
    .B(\game.ballX[8] ),
    .Y(_0349_));
 sky130_fd_sc_hd__a21oi_1 _0800_ (.A1(\game.ballX[7] ),
    .A2(_0346_),
    .B1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__or2_1 _0801_ (.A(_0064_),
    .B(\game.ballX[0] ),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _0802_ (.A(_0064_),
    .B(\game.ballX[0] ),
    .Y(_0352_));
 sky130_fd_sc_hd__or2_1 _0803_ (.A(_0065_),
    .B(\game.ballX[1] ),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _0804_ (.A(_0065_),
    .B(\game.ballX[1] ),
    .Y(_0354_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0353_),
    .B2(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__xnor2_1 _0806_ (.A(_0066_),
    .B(\game.ballX[3] ),
    .Y(_0356_));
 sky130_fd_sc_hd__xnor2_1 _0807_ (.A(\game.h[3] ),
    .B(\game.ballX[2] ),
    .Y(_0357_));
 sky130_fd_sc_hd__nand3_1 _0808_ (.A(\game.ballX[3] ),
    .B(_0292_),
    .C(\game.ballX[5] ),
    .Y(_0358_));
 sky130_fd_sc_hd__xor2_2 _0809_ (.A(\game.h[7] ),
    .B(\game.ballX[6] ),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_1 _0810_ (.A(\game.ballX[3] ),
    .B(_0292_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _0811_ (.A(_0130_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__a22oi_1 _0812_ (.A1(_0358_),
    .A2(_0359_),
    .B1(_0361_),
    .B2(_0063_),
    .Y(_0362_));
 sky130_fd_sc_hd__or4bb_1 _0813_ (.A(_0355_),
    .B(_0356_),
    .C_N(_0357_),
    .D_N(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__xnor2_1 _0814_ (.A(\game.h[6] ),
    .B(\game.ballX[5] ),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_1 _0815_ (.A(_0130_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__a21o_1 _0816_ (.A1(\game.ballX[3] ),
    .A2(_0292_),
    .B1(_0364_),
    .X(_0366_));
 sky130_fd_sc_hd__o221a_1 _0817_ (.A1(_0358_),
    .A2(_0359_),
    .B1(_0365_),
    .B2(_0063_),
    .C1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__or4b_1 _0818_ (.A(_0348_),
    .B(_0350_),
    .C(_0363_),
    .D_N(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(_0359_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_1 _0820_ (.A(_0063_),
    .B(_0292_),
    .Y(_0370_));
 sky130_fd_sc_hd__and4_1 _0821_ (.A(_0347_),
    .B(_0356_),
    .C(_0357_),
    .D(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__and4b_1 _0822_ (.A_N(_0355_),
    .B(_0364_),
    .C(_0369_),
    .D(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__a31o_1 _0823_ (.A1(\game.inBallX ),
    .A2(\game.ballX[7] ),
    .A3(_0346_),
    .B1(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__a22o_1 _0824_ (.A1(\game.inBallX ),
    .A2(_0368_),
    .B1(_0373_),
    .B2(_0349_),
    .X(_0374_));
 sky130_fd_sc_hd__a211o_1 _0825_ (.A1(_0292_),
    .A2(\game.ballX[5] ),
    .B1(\game.ballX[6] ),
    .C1(\game.ballX[7] ),
    .X(_0375_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(\game.ballX[8] ),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__and3_1 _0827_ (.A(_0138_),
    .B(_0374_),
    .C(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0828_ (.A(_0377_),
    .X(_0032_));
 sky130_fd_sc_hd__o21ai_1 _0829_ (.A1(_0059_),
    .A2(_0078_),
    .B1(net15),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(\game.inBallY ),
    .Y(_0379_));
 sky130_fd_sc_hd__o21ai_1 _0831_ (.A1(_0379_),
    .A2(_0081_),
    .B1(_0244_),
    .Y(_0380_));
 sky130_fd_sc_hd__a21o_1 _0832_ (.A1(_0378_),
    .A2(_0380_),
    .B1(_0209_),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(\game.inBallX ),
    .Y(_0381_));
 sky130_fd_sc_hd__o21a_1 _0834_ (.A1(_0381_),
    .A2(_0080_),
    .B1(_0295_),
    .X(_0382_));
 sky130_fd_sc_hd__or3_1 _0835_ (.A(_0209_),
    .B(_0343_),
    .C(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(_0383_),
    .X(_0034_));
 sky130_fd_sc_hd__and3_1 _0837_ (.A(\game.ballY[3] ),
    .B(\game.ballY[4] ),
    .C(\game.ballY[5] ),
    .X(_0384_));
 sky130_fd_sc_hd__nand3_1 _0838_ (.A(\game.ballY[6] ),
    .B(\game.ballY[7] ),
    .C(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__xor2_1 _0839_ (.A(\game.v[7] ),
    .B(\game.ballY[6] ),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _0840_ (.A(_0386_),
    .B(_0384_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(_0386_),
    .B(_0384_),
    .Y(_0388_));
 sky130_fd_sc_hd__xnor2_1 _0842_ (.A(\game.v[8] ),
    .B(\game.ballY[7] ),
    .Y(_0389_));
 sky130_fd_sc_hd__and3_1 _0843_ (.A(\game.ballY[6] ),
    .B(_0389_),
    .C(_0384_),
    .X(_0390_));
 sky130_fd_sc_hd__a221o_1 _0844_ (.A1(_0059_),
    .A2(_0385_),
    .B1(_0387_),
    .B2(_0388_),
    .C1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__a21oi_1 _0845_ (.A1(\game.ballY[6] ),
    .A2(_0384_),
    .B1(_0389_),
    .Y(_0392_));
 sky130_fd_sc_hd__xnor2_1 _0846_ (.A(_0084_),
    .B(\game.ballY[4] ),
    .Y(_0393_));
 sky130_fd_sc_hd__xnor2_1 _0847_ (.A(\game.v[6] ),
    .B(\game.ballY[5] ),
    .Y(_0394_));
 sky130_fd_sc_hd__o21ai_1 _0848_ (.A1(\game.ballY[3] ),
    .A2(_0393_),
    .B1(_0142_),
    .Y(_0395_));
 sky130_fd_sc_hd__a221o_1 _0849_ (.A1(\game.ballY[3] ),
    .A2(_0393_),
    .B1(_0394_),
    .B2(_0133_),
    .C1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(_0059_),
    .B(_0385_),
    .Y(_0397_));
 sky130_fd_sc_hd__or2_1 _0851_ (.A(\game.v[2] ),
    .B(\game.ballY[1] ),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _0852_ (.A(\game.v[2] ),
    .B(\game.ballY[1] ),
    .Y(_0399_));
 sky130_fd_sc_hd__xor2_1 _0853_ (.A(\game.v[1] ),
    .B(\game.ballY[0] ),
    .X(_0400_));
 sky130_fd_sc_hd__a21oi_1 _0854_ (.A1(_0398_),
    .A2(_0399_),
    .B1(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_1 _0855_ (.A(\game.v[3] ),
    .B(\game.ballY[2] ),
    .Y(_0402_));
 sky130_fd_sc_hd__xor2_1 _0856_ (.A(\game.v[4] ),
    .B(\game.ballY[3] ),
    .X(_0403_));
 sky130_fd_sc_hd__and3_1 _0857_ (.A(\game.inBallY ),
    .B(_0402_),
    .C(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__o211a_1 _0858_ (.A1(_0133_),
    .A2(_0394_),
    .B1(_0401_),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__or4b_1 _0859_ (.A(_0392_),
    .B(_0396_),
    .C(_0397_),
    .D_N(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__and4b_1 _0860_ (.A_N(_0386_),
    .B(_0393_),
    .C(_0394_),
    .D(_0402_),
    .X(_0407_));
 sky130_fd_sc_hd__and3b_1 _0861_ (.A_N(_0403_),
    .B(_0401_),
    .C(_0389_),
    .X(_0408_));
 sky130_fd_sc_hd__a31o_1 _0862_ (.A1(_0142_),
    .A2(_0407_),
    .A3(_0408_),
    .B1(\game.inBallY ),
    .X(_0409_));
 sky130_fd_sc_hd__o211a_1 _0863_ (.A1(_0391_),
    .A2(_0406_),
    .B1(_0161_),
    .C1(_0409_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_2 _0864_ (.A(_0208_),
    .B(_0142_),
    .Y(_0410_));
 sky130_fd_sc_hd__and2b_1 _0865_ (.A_N(_0062_),
    .B(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0866_ (.A(_0411_),
    .X(_0036_));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(_0064_),
    .B(_0062_),
    .Y(_0412_));
 sky130_fd_sc_hd__or2_1 _0868_ (.A(_0064_),
    .B(_0062_),
    .X(_0413_));
 sky130_fd_sc_hd__and3_1 _0869_ (.A(_0412_),
    .B(_0410_),
    .C(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _0870_ (.A(_0414_),
    .X(_0037_));
 sky130_fd_sc_hd__nand3_1 _0871_ (.A(_0064_),
    .B(_0062_),
    .C(_0065_),
    .Y(_0415_));
 sky130_fd_sc_hd__a21o_1 _0872_ (.A1(_0064_),
    .A2(_0062_),
    .B1(_0065_),
    .X(_0416_));
 sky130_fd_sc_hd__and3_1 _0873_ (.A(_0138_),
    .B(_0415_),
    .C(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0417_),
    .X(_0038_));
 sky130_fd_sc_hd__a31o_1 _0875_ (.A1(_0064_),
    .A2(_0062_),
    .A3(_0065_),
    .B1(\game.h[3] ),
    .X(_0418_));
 sky130_fd_sc_hd__and3b_1 _0876_ (.A_N(_0140_),
    .B(_0418_),
    .C(net1),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _0877_ (.A(_0419_),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _0878_ (.A(_0066_),
    .B(_0140_),
    .X(_0420_));
 sky130_fd_sc_hd__o21ai_1 _0879_ (.A1(_0066_),
    .A2(_0140_),
    .B1(_0410_),
    .Y(_0421_));
 sky130_fd_sc_hd__nor2_1 _0880_ (.A(_0420_),
    .B(_0421_),
    .Y(_0040_));
 sky130_fd_sc_hd__o21ai_1 _0881_ (.A1(_0063_),
    .A2(_0420_),
    .B1(_0410_),
    .Y(_0422_));
 sky130_fd_sc_hd__a21oi_1 _0882_ (.A1(_0063_),
    .A2(_0420_),
    .B1(_0422_),
    .Y(_0041_));
 sky130_fd_sc_hd__and3_1 _0883_ (.A(_0066_),
    .B(_0079_),
    .C(_0140_),
    .X(_0423_));
 sky130_fd_sc_hd__a31o_1 _0884_ (.A1(_0063_),
    .A2(_0066_),
    .A3(_0140_),
    .B1(\game.h[6] ),
    .X(_0424_));
 sky130_fd_sc_hd__and3b_1 _0885_ (.A_N(_0423_),
    .B(_0410_),
    .C(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _0886_ (.A(_0425_),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _0887_ (.A(\game.h[7] ),
    .B(_0423_),
    .X(_0426_));
 sky130_fd_sc_hd__o21ai_1 _0888_ (.A1(net22),
    .A2(_0423_),
    .B1(_0410_),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_1 _0889_ (.A(_0426_),
    .B(_0427_),
    .Y(_0043_));
 sky130_fd_sc_hd__and3_1 _0890_ (.A(\game.h[7] ),
    .B(\game.h[8] ),
    .C(_0423_),
    .X(_0428_));
 sky130_fd_sc_hd__or2_1 _0891_ (.A(\game.h[8] ),
    .B(_0426_),
    .X(_0429_));
 sky130_fd_sc_hd__and3b_1 _0892_ (.A_N(_0428_),
    .B(_0410_),
    .C(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _0893_ (.A(_0430_),
    .X(_0044_));
 sky130_fd_sc_hd__o21ai_1 _0894_ (.A1(net11),
    .A2(_0428_),
    .B1(_0410_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21oi_1 _0895_ (.A1(net11),
    .A2(_0428_),
    .B1(_0431_),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2_1 _0896_ (.A(\game.paddle[7] ),
    .B(\game.paddle[6] ),
    .Y(_0432_));
 sky130_fd_sc_hd__xnor2_1 _0897_ (.A(_0432_),
    .B(_0340_),
    .Y(_0433_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(_0337_),
    .A1(_0338_),
    .S(_0339_),
    .X(_0434_));
 sky130_fd_sc_hd__and3_1 _0899_ (.A(\game.paddle[7] ),
    .B(\game.paddle[6] ),
    .C(\game.paddle[8] ),
    .X(_0435_));
 sky130_fd_sc_hd__xor2_1 _0900_ (.A(_0059_),
    .B(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__o41a_1 _0901_ (.A1(_0336_),
    .A2(_0433_),
    .A3(_0434_),
    .A4(_0436_),
    .B1(net16),
    .X(_0437_));
 sky130_fd_sc_hd__o21a_1 _0902_ (.A1(_0342_),
    .A2(_0437_),
    .B1(_0161_),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _0903_ (.A(\game.v[0] ),
    .B(_0142_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_1 _0904_ (.A(_0208_),
    .B(net6),
    .Y(_0439_));
 sky130_fd_sc_hd__o21ai_1 _0905_ (.A1(net21),
    .A2(_0142_),
    .B1(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _0906_ (.A(_0438_),
    .B(_0440_),
    .Y(_0047_));
 sky130_fd_sc_hd__and3_1 _0907_ (.A(\game.v[1] ),
    .B(\game.v[0] ),
    .C(_0142_),
    .X(_0441_));
 sky130_fd_sc_hd__or2_1 _0908_ (.A(\game.v[1] ),
    .B(_0438_),
    .X(_0442_));
 sky130_fd_sc_hd__and3b_1 _0909_ (.A_N(_0441_),
    .B(_0138_),
    .C(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0910_ (.A(_0443_),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(\game.v[2] ),
    .B(_0441_),
    .X(_0444_));
 sky130_fd_sc_hd__or2_1 _0912_ (.A(\game.v[2] ),
    .B(_0441_),
    .X(_0445_));
 sky130_fd_sc_hd__and3b_1 _0913_ (.A_N(_0444_),
    .B(_0439_),
    .C(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0914_ (.A(_0446_),
    .X(_0049_));
 sky130_fd_sc_hd__and3_1 _0915_ (.A(\game.v[3] ),
    .B(\game.v[2] ),
    .C(_0441_),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _0916_ (.A(\game.v[3] ),
    .B(_0444_),
    .X(_0448_));
 sky130_fd_sc_hd__and3b_1 _0917_ (.A_N(_0447_),
    .B(_0439_),
    .C(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _0918_ (.A(_0449_),
    .X(_0050_));
 sky130_fd_sc_hd__and3_1 _0919_ (.A(\game.v[4] ),
    .B(\game.v[3] ),
    .C(_0444_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(\game.v[4] ),
    .B(_0447_),
    .X(_0451_));
 sky130_fd_sc_hd__and3b_1 _0921_ (.A_N(_0450_),
    .B(_0138_),
    .C(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0922_ (.A(_0452_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _0923_ (.A(_0084_),
    .B(_0450_),
    .X(_0453_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(_0084_),
    .B(_0450_),
    .X(_0454_));
 sky130_fd_sc_hd__and3b_1 _0925_ (.A_N(_0453_),
    .B(net1),
    .C(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0926_ (.A(_0455_),
    .X(_0052_));
 sky130_fd_sc_hd__a31o_1 _0927_ (.A1(\game.v[6] ),
    .A2(_0084_),
    .A3(_0450_),
    .B1(_0209_),
    .X(_0456_));
 sky130_fd_sc_hd__o21ba_1 _0928_ (.A1(net20),
    .A2(_0453_),
    .B1_N(_0456_),
    .X(_0053_));
 sky130_fd_sc_hd__and3_1 _0929_ (.A(\game.v[7] ),
    .B(\game.v[6] ),
    .C(_0453_),
    .X(_0457_));
 sky130_fd_sc_hd__a31o_1 _0930_ (.A1(\game.v[6] ),
    .A2(_0084_),
    .A3(_0450_),
    .B1(\game.v[7] ),
    .X(_0458_));
 sky130_fd_sc_hd__and3b_1 _0931_ (.A_N(_0457_),
    .B(net1),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _0932_ (.A(_0459_),
    .X(_0054_));
 sky130_fd_sc_hd__and3_1 _0933_ (.A(_0084_),
    .B(_0078_),
    .C(_0450_),
    .X(_0460_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__o211a_1 _0935_ (.A1(net18),
    .A2(_0457_),
    .B1(_0461_),
    .C1(_0161_),
    .X(_0055_));
 sky130_fd_sc_hd__o21ai_1 _0936_ (.A1(_0059_),
    .A2(_0460_),
    .B1(_0439_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21oi_1 _0937_ (.A1(_0059_),
    .A2(_0460_),
    .B1(_0462_),
    .Y(_0056_));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0000_),
    .Q(\game.offset[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0001_),
    .Q(\game.offset[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0940_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0002_),
    .Q(\game.offset[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0003_),
    .Q(\game.offset[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0004_),
    .Q(\game.offset[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0005_),
    .Q(\game.paddle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0944_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0006_),
    .Q(\game.paddle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0945_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0007_),
    .Q(\game.paddle[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0946_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0008_),
    .Q(\game.paddle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0947_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0009_),
    .Q(\game.paddle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _0948_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0010_),
    .Q(\game.paddle[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0949_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0011_),
    .Q(\game.paddle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0950_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0012_),
    .Q(\game.paddle[7] ));
 sky130_fd_sc_hd__dfxtp_2 _0951_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0013_),
    .Q(\game.paddle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_3_3__leaf_clk),
    .D(\game.red ),
    .Q(qr));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_3_3__leaf_clk),
    .D(\game.green ),
    .Q(qg));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_3_6__leaf_clk),
    .D(\game.blue ),
    .Q(qb));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_3_7__leaf_clk),
    .D(net10),
    .Q(\game.pause_n ));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_3_7__leaf_clk),
    .D(\pause.d ),
    .Q(\pause.dff1 ));
 sky130_fd_sc_hd__dfxtp_2 _0957_ (.CLK(clknet_3_7__leaf_clk),
    .D(net9),
    .Q(\game.new_game_n ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_3_7__leaf_clk),
    .D(\new_game.d ),
    .Q(\new_game.dff1 ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_3_7__leaf_clk),
    .D(net8),
    .Q(\down_key.dff2 ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_3_7__leaf_clk),
    .D(\down_key.d ),
    .Q(\down_key.dff1 ));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_3_7__leaf_clk),
    .D(net7),
    .Q(\game.up_key_n ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_3_6__leaf_clk),
    .D(\up_key.d ),
    .Q(\up_key.dff1 ));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0014_),
    .Q(\game.ballY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0964_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0015_),
    .Q(\game.ballY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0016_),
    .Q(\game.ballY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0966_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0017_),
    .Q(\game.ballY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0018_),
    .Q(\game.ballY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0019_),
    .Q(\game.ballY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0969_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0020_),
    .Q(\game.ballY[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0970_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0021_),
    .Q(\game.ballY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0022_),
    .Q(\game.ballX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0023_),
    .Q(\game.ballX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0024_),
    .Q(\game.ballX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0974_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0025_),
    .Q(\game.ballX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0026_),
    .Q(\game.ballX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _0976_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0027_),
    .Q(\game.ballX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0977_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0028_),
    .Q(\game.ballX[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0978_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0029_),
    .Q(\game.ballX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0030_),
    .Q(\game.ballX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0031_),
    .Q(\game.hit ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0032_),
    .Q(\game.inBallX ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0033_),
    .Q(\game.ballDirY ));
 sky130_fd_sc_hd__dfxtp_2 _0983_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0034_),
    .Q(\game.ballDirX ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0035_),
    .Q(\game.inBallY ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0036_),
    .Q(\game.h[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0037_),
    .Q(\game.h[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0038_),
    .Q(\game.h[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0988_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0039_),
    .Q(\game.h[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0040_),
    .Q(\game.h[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0041_),
    .Q(\game.h[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0042_),
    .Q(\game.h[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0992_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0043_),
    .Q(\game.h[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0044_),
    .Q(\game.h[8] ));
 sky130_fd_sc_hd__dfxtp_2 _0994_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0045_),
    .Q(\game.h[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0046_),
    .Q(\game.inPaddle ));
 sky130_fd_sc_hd__dfxtp_2 _0996_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0047_),
    .Q(\game.v[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0997_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0048_),
    .Q(\game.v[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0998_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0049_),
    .Q(\game.v[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0999_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0050_),
    .Q(\game.v[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1000_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0051_),
    .Q(\game.v[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0052_),
    .Q(\game.v[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1002_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0053_),
    .Q(\game.v[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0054_),
    .Q(\game.v[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1004_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0055_),
    .Q(\game.v[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0056_),
    .Q(\game.v[9] ));
 sky130_fd_sc_hd__clkbuf_4 _1006_ (.A(qb),
    .X(uo_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _1007_ (.A(qg),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _1008_ (.A(qr),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _1009_ (.A(\game.hsync ),
    .X(uo_out[3]));
 sky130_fd_sc_hd__clkbuf_4 _1010_ (.A(\game.vsync ),
    .X(uo_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _1011_ (.A(\game.speaker ),
    .X(uo_out[5]));
 sky130_fd_sc_hd__clkbuf_4 _1012_ (.A(\game.col0 ),
    .X(uo_out[6]));
 sky130_fd_sc_hd__clkbuf_4 _1013_ (.A(\game.row0 ),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\up_key.dff1 ),
    .X(net7));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\game.inPaddle ),
    .X(net16));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\game.paddle[6] ),
    .X(net17));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\game.v[8] ),
    .X(net18));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\game.paddle[0] ),
    .X(net19));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\game.v[6] ),
    .X(net20));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\game.v[0] ),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\game.h[7] ),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\game.inBallX ),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\down_key.dff1 ),
    .X(net8));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\new_game.dff1 ),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\pause.dff1 ),
    .X(net10));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\game.h[9] ),
    .X(net11));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\game.offset[4] ),
    .X(net12));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\game.ballY[7] ),
    .X(net13));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\game.ballX[6] ),
    .X(net14));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\game.inBallY ),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 max_cap6 (.A(_0152_),
    .X(net6));
endmodule

