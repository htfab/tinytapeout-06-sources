magic
tech sky130A
magscale 1 2
timestamp 1713144495
<< pwell >>
rect 5300 480 5330 690
rect 2080 -1100 2240 -1020
rect 2340 -1100 2500 -1020
<< locali >>
rect 1460 1880 5640 2100
rect 1460 1280 1860 1880
rect 2160 1640 2300 1880
rect 2680 1640 2820 1880
rect 3100 1280 3660 1880
rect 3960 1640 4100 1880
rect 4460 1640 4600 1880
rect 4900 1280 5640 1880
rect 1460 1020 5640 1280
rect 1520 760 5650 900
rect 1520 700 4080 760
rect 5290 740 5650 760
rect 5300 720 5650 740
rect 1520 -1120 1660 700
rect 2920 614 4060 700
rect 2920 -24 3216 614
rect 3694 -24 4060 614
rect 2920 -270 4060 -24
rect 2920 -880 3120 -270
rect 3840 -280 4060 -270
rect 3440 -880 3540 -420
rect 3860 -880 4060 -280
rect 5300 -680 5420 720
rect 2920 -1120 4060 -880
rect 5310 -1120 5420 -680
rect 1510 -1200 5420 -1120
rect 5550 -1200 5650 720
rect 1510 -1240 5650 -1200
rect 1510 -1370 1720 -1240
rect 5280 -1370 5650 -1240
rect 1510 -1420 5650 -1370
rect 1510 -1430 5390 -1420
<< viali >>
rect 3216 -24 3694 614
rect 5420 -1200 5550 720
rect 1720 -1370 5280 -1240
<< metal1 >>
rect 1460 1840 5640 2100
rect 1520 1820 3080 1840
rect 3640 1820 5640 1840
rect 2160 1640 2300 1820
rect 2680 1640 2820 1820
rect 3960 1640 4100 1820
rect 4460 1640 4600 1820
rect 2980 1600 3320 1620
rect 2980 1580 3100 1600
rect 1920 1430 3100 1580
rect 3300 1430 3320 1600
rect 1920 1420 3320 1430
rect 3420 1600 3800 1620
rect 3420 1440 3440 1600
rect 3660 1440 4860 1600
rect 3420 1420 4860 1440
rect 1460 1260 4940 1380
rect 3400 970 3570 976
rect 1445 800 3400 970
rect 3400 794 3570 800
rect 3990 760 5650 900
rect 1520 700 2940 750
rect 1520 -1120 1660 700
rect 1720 550 1840 620
rect 1720 -50 1740 550
rect 1800 -50 1840 550
rect 1720 -70 1840 -50
rect 2220 580 2340 630
rect 2220 -20 2250 580
rect 2310 -20 2340 580
rect 2220 -60 2340 -20
rect 2720 570 2840 630
rect 2720 -30 2750 570
rect 2810 -30 2840 570
rect 2720 -60 2840 -30
rect 2908 620 2940 700
rect 4010 700 4080 760
rect 5290 740 5650 760
rect 5300 720 5650 740
rect 4010 630 4054 700
rect 3970 620 4054 630
rect 2908 614 4054 620
rect 2908 -24 3216 614
rect 3694 -24 4054 614
rect 2908 -90 4054 -24
rect 4110 550 4230 600
rect 4110 -50 4130 550
rect 4190 -50 4230 550
rect 4110 -90 4230 -50
rect 4620 560 4740 600
rect 4620 -40 4650 560
rect 4710 -40 4740 560
rect 4620 -90 4740 -40
rect 5130 550 5250 600
rect 5130 -50 5150 550
rect 5210 -50 5250 550
rect 5130 -90 5250 -50
rect 2908 -140 3110 -90
rect 2900 -270 3110 -140
rect 3860 -120 4054 -90
rect 3360 -180 3610 -150
rect 3360 -240 3430 -180
rect 3530 -240 3610 -180
rect 3360 -270 3610 -240
rect 3860 -270 4060 -120
rect 1960 -440 2080 -420
rect 1960 -700 2000 -440
rect 2060 -700 2080 -440
rect 1960 -720 2080 -700
rect 2480 -440 2600 -420
rect 2480 -700 2500 -440
rect 2560 -700 2600 -440
rect 2480 -720 2600 -700
rect 2900 -880 3120 -270
rect 3430 -300 3530 -270
rect 3240 -380 3760 -300
rect 3180 -440 3280 -420
rect 3180 -700 3200 -440
rect 3260 -700 3280 -440
rect 3180 -720 3280 -700
rect 3440 -880 3540 -420
rect 3700 -440 3800 -420
rect 3760 -700 3800 -440
rect 3700 -720 3800 -700
rect 3840 -880 4060 -270
rect 4380 -440 4480 -420
rect 4440 -700 4480 -440
rect 4380 -720 4480 -700
rect 4900 -440 5000 -420
rect 4960 -700 5000 -440
rect 5300 -680 5420 720
rect 4900 -720 5000 -700
rect 1780 -1100 1820 -1020
rect 1980 -1100 2080 -1020
rect 2240 -1100 2340 -1020
rect 2500 -1100 2600 -1020
rect 2760 -1100 2800 -1020
rect 2900 -1120 4060 -880
rect 4160 -1100 4220 -1020
rect 4380 -1100 4480 -1020
rect 4640 -1100 4740 -1020
rect 4900 -1100 5000 -1020
rect 5160 -1100 5220 -1020
rect 5310 -1120 5420 -680
rect 1520 -1140 1740 -1120
rect 2840 -1140 4080 -1120
rect 4132 -1140 5234 -1130
rect 5280 -1140 5420 -1120
rect 1510 -1200 5420 -1140
rect 5550 -1200 5650 720
rect 1510 -1240 5650 -1200
rect 1510 -1370 1720 -1240
rect 5280 -1370 5650 -1240
rect 1510 -1420 5650 -1370
rect 1510 -1430 5380 -1420
<< via1 >>
rect 3100 1430 3300 1600
rect 3440 1440 3660 1600
rect 3400 800 3570 970
rect 1740 -50 1800 550
rect 2250 -20 2310 580
rect 2750 -30 2810 570
rect 4130 -50 4190 550
rect 4650 -40 4710 560
rect 5150 -50 5210 550
rect 3430 -240 3530 -180
rect 2000 -700 2060 -440
rect 2500 -700 2560 -440
rect 3200 -700 3260 -440
rect 3700 -700 3760 -440
rect 4380 -700 4440 -440
rect 4900 -700 4960 -440
rect 1820 -1100 1980 -1020
rect 2080 -1100 2240 -1020
rect 2340 -1100 2500 -1020
rect 2600 -1100 2760 -1020
rect 4220 -1100 4380 -1020
rect 4480 -1100 4640 -1020
rect 4740 -1100 4900 -1020
rect 5000 -1100 5160 -1020
<< metal2 >>
rect 3100 1660 3340 2100
rect 3080 1600 3340 1660
rect 3080 1430 3100 1600
rect 3300 1430 3340 1600
rect 3080 1420 3340 1430
rect 3420 1660 3660 2100
rect 3420 1600 3680 1660
rect 3420 1440 3440 1600
rect 3660 1440 3680 1600
rect 3420 1420 3680 1440
rect 1720 580 2900 610
rect 1720 550 2250 580
rect 1720 -50 1740 550
rect 1800 -20 2250 550
rect 2310 570 2900 580
rect 2310 -20 2750 570
rect 1800 -30 2750 -20
rect 2810 349 2900 570
rect 3102 349 3319 1420
rect 3440 1190 3660 1420
rect 3440 1030 3970 1190
rect 3394 800 3400 970
rect 3570 800 3576 970
rect 3740 940 3970 1030
rect 2810 132 3319 349
rect 2810 -30 2900 132
rect 1800 -50 2900 -30
rect 1720 -160 2900 -50
rect 3400 -180 3570 800
rect 3750 350 3970 940
rect 4090 560 5270 600
rect 4090 550 4650 560
rect 4090 350 4130 550
rect 3750 130 4130 350
rect 4090 -50 4130 130
rect 4190 -40 4650 550
rect 4710 550 5270 560
rect 4710 -40 5150 550
rect 4190 -50 5150 -40
rect 5210 -50 5270 550
rect 4090 -170 5270 -50
rect 3400 -240 3430 -180
rect 3530 -240 3570 -180
rect 3400 -260 3570 -240
rect 1960 -440 5020 -420
rect 1960 -700 2000 -440
rect 2060 -700 2500 -440
rect 2560 -700 3200 -440
rect 3260 -700 3700 -440
rect 3760 -700 4380 -440
rect 4440 -700 4900 -440
rect 4960 -700 5020 -440
rect 1960 -720 5020 -700
rect 3100 -1020 3320 -960
rect 1780 -1100 1820 -1020
rect 1980 -1100 2080 -1020
rect 2240 -1100 2340 -1020
rect 2500 -1100 2600 -1020
rect 2760 -1100 3320 -1020
rect 3100 -1420 3320 -1100
rect 3600 -1020 3820 -960
rect 3600 -1100 4220 -1020
rect 4380 -1100 4480 -1020
rect 4640 -1100 4740 -1020
rect 4900 -1100 5000 -1020
rect 5160 -1100 5220 -1020
rect 3600 -1420 3820 -1100
use sky130_fd_pr__nfet_01v8_5WCAAQ  sky130_fd_pr__nfet_01v8_5WCAAQ_0
timestamp 1713067979
transform -1 0 2283 0 1 -221
box -683 -979 683 979
use sky130_fd_pr__nfet_01v8_JL39Q5  sky130_fd_pr__nfet_01v8_JL39Q5_0
timestamp 1713142989
transform 1 0 3485 0 1 -581
box -425 -379 425 379
use sky130_fd_pr__nfet_01v8_MM2THM  sky130_fd_pr__nfet_01v8_MM2THM_0
timestamp 1713067979
transform 1 0 4683 0 1 -190
box -683 -1010 683 1010
use sky130_fd_pr__pfet_01v8_D6KM8H  sky130_fd_pr__pfet_01v8_D6KM8H_0
timestamp 1713067979
transform 1 0 2483 0 1 1584
box -683 -384 683 384
use sky130_fd_pr__pfet_01v8_D6KM8H  sky130_fd_pr__pfet_01v8_D6KM8H_1
timestamp 1713067979
transform 1 0 4283 0 1 1584
box -683 -384 683 384
<< labels >>
flabel metal2 3140 -1100 3240 -1020 0 FreeSans 1600 270 0 0 VIN_N
port 1 nsew
flabel metal2 3680 -1100 3780 -1020 0 FreeSans 1600 270 0 0 VIN
port 0 nsew
flabel metal1 1520 1820 1820 1980 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
flabel metal1 1520 -1260 1680 -1140 0 FreeSans 1600 0 0 0 VSS
port 7 nsew
flabel metal1 1460 1260 1580 1380 0 FreeSans 1600 0 0 0 VPBIAS
port 8 nsew
flabel metal1 1445 800 1615 970 0 FreeSans 1600 0 0 0 VNBIAS
port 5 nsew
flabel metal2 3100 1860 3340 2100 0 FreeSans 1600 270 0 0 VOUT
port 2 nsew
flabel metal2 3420 1860 3660 2100 0 FreeSans 1600 270 0 0 VOUT_N
port 3 nsew
<< end >>
