magic
tech sky130A
timestamp 1713125316
<< metal1 >>
rect 5358 2758 13797 2773
rect 5358 2683 5369 2758
rect 5526 2683 13797 2758
rect 5358 2671 13797 2683
rect 14325 2195 15715 2208
rect 14325 2119 15592 2195
rect 15705 2119 15715 2195
rect 14325 2108 15715 2119
rect 9032 1959 10379 1973
rect 9032 1842 9046 1959
rect 9172 1873 10379 1959
rect 9172 1842 9185 1873
rect 14329 1859 15419 1959
rect 9032 1829 9185 1842
rect 14331 1640 14902 1740
rect 9538 1281 13796 1300
rect 9538 1215 9555 1281
rect 9681 1215 13796 1281
rect 9538 1198 13796 1215
rect 14826 812 14902 1640
rect 11239 803 14902 812
rect 11239 741 11253 803
rect 11397 741 14902 803
rect 11239 731 14902 741
rect 15328 524 15419 1859
rect 13448 513 15419 524
rect 13448 459 13460 513
rect 13551 459 15419 513
rect 13448 446 15419 459
<< via1 >>
rect 5369 2683 5526 2758
rect 15592 2119 15705 2195
rect 9046 1842 9172 1959
rect 9555 1215 9681 1281
rect 11253 741 11397 803
rect 13460 459 13551 513
<< metal2 >>
rect 5357 2758 5539 2774
rect 5357 2683 5369 2758
rect 5526 2683 5539 2758
rect 5357 2670 5539 2683
rect 15577 2195 15716 2208
rect 15577 2119 15592 2195
rect 15705 2119 15716 2195
rect 15577 2108 15716 2119
rect 9032 1959 9186 1974
rect 9032 1842 9046 1959
rect 9172 1842 9186 1959
rect 9032 1828 9186 1842
rect 581 1300 5627 1304
rect 581 1291 9699 1300
rect 581 1207 592 1291
rect 729 1281 9699 1291
rect 729 1215 9555 1281
rect 9681 1215 9699 1281
rect 729 1207 9699 1215
rect 581 1197 9699 1207
rect 5546 1196 9699 1197
rect 11239 803 11408 812
rect 11239 741 11253 803
rect 11397 741 11408 803
rect 11239 731 11408 741
rect 13448 513 13561 524
rect 13448 459 13460 513
rect 13551 459 13561 513
rect 13448 446 13561 459
<< via2 >>
rect 5369 2683 5526 2758
rect 15592 2119 15705 2195
rect 9046 1842 9172 1959
rect 592 1207 729 1291
rect 11253 741 11397 803
rect 13460 459 13551 513
<< metal3 >>
rect 5357 2758 5539 2774
rect 5357 2683 5369 2758
rect 5526 2683 5539 2758
rect 5357 2670 5539 2683
rect 15577 2195 15716 2208
rect 15577 2119 15592 2195
rect 15705 2119 15716 2195
rect 15577 2108 15716 2119
rect 9032 1959 9186 1974
rect 9032 1842 9046 1959
rect 9172 1842 9186 1959
rect 9032 1828 9186 1842
rect 581 1291 739 1304
rect 581 1207 592 1291
rect 729 1207 739 1291
rect 581 1197 739 1207
rect 11239 803 11408 812
rect 11239 741 11253 803
rect 11397 741 11408 803
rect 11239 731 11408 741
rect 13448 513 13561 524
rect 13448 459 13460 513
rect 13551 459 13561 513
rect 13448 446 13561 459
<< via3 >>
rect 5369 2683 5526 2758
rect 15592 2119 15705 2195
rect 9046 1842 9172 1959
rect 592 1207 729 1291
rect 11253 741 11397 803
rect 13460 459 13551 513
<< metal4 >>
rect 399 22412 429 22576
rect 767 22412 797 22576
rect 1135 22412 1165 22576
rect 1503 22412 1533 22576
rect 1871 22412 1901 22576
rect 2239 22412 2269 22576
rect 2607 22412 2637 22576
rect 2975 22412 3005 22576
rect 3343 22412 3373 22576
rect 3711 22412 3741 22576
rect 4079 22412 4109 22576
rect 4447 22412 4477 22576
rect 4815 22412 4845 22576
rect 5183 22412 5213 22576
rect 5551 22412 5581 22576
rect 5919 22412 5949 22576
rect 6287 22412 6317 22576
rect 6655 22412 6685 22576
rect 7023 22412 7053 22576
rect 7391 22412 7421 22576
rect 7759 22412 7789 22576
rect 8127 22412 8157 22576
rect 8495 22412 8525 22576
rect 8863 22412 8893 22576
rect 9231 22451 9261 22576
rect 9599 22451 9629 22576
rect 9967 22451 9997 22576
rect 10335 22451 10365 22576
rect 10703 22451 10733 22576
rect 11071 22451 11101 22576
rect 11439 22451 11469 22576
rect 11807 22451 11837 22576
rect 12175 22451 12205 22576
rect 12543 22451 12573 22576
rect 12911 22451 12941 22576
rect 13279 22451 13309 22576
rect 13647 22451 13677 22576
rect 14015 22451 14045 22576
rect 14383 22451 14413 22576
rect 14751 22451 14781 22576
rect 15119 22451 15149 22576
rect 15487 22451 15517 22576
rect 15855 22451 15885 22576
rect 399 22309 8894 22412
rect 100 1304 250 22076
rect 4900 2774 5050 22309
rect 4900 2758 5539 2774
rect 4900 2683 5369 2758
rect 5526 2683 5539 2758
rect 4900 2671 5539 2683
rect 4900 1436 5050 2671
rect 15577 2195 15716 2208
rect 15577 2119 15592 2195
rect 15705 2119 15716 2195
rect 15577 2108 15716 2119
rect 9032 1959 9185 1973
rect 9032 1842 9046 1959
rect 9172 1842 9185 1959
rect 9032 1829 9185 1842
rect 100 1291 739 1304
rect 100 1207 592 1291
rect 729 1207 739 1291
rect 100 1197 739 1207
rect 100 1196 251 1197
rect 100 500 250 1196
rect 4900 1063 5049 1436
rect 9032 1204 9092 1829
rect 9031 1082 9092 1204
rect 4900 500 5050 1063
rect 200 0 260 100
rect 2408 0 2468 100
rect 4616 0 4676 100
rect 6824 0 6884 100
rect 9032 0 9092 1082
rect 11239 803 11408 812
rect 11239 741 11253 803
rect 11397 741 11408 803
rect 11239 731 11408 741
rect 11239 89 11301 731
rect 13448 513 13561 524
rect 13448 459 13460 513
rect 13551 459 13561 513
rect 13448 446 13561 459
rect 11240 0 11300 89
rect 13448 0 13508 446
rect 15655 100 15715 2108
rect 15655 88 15716 100
rect 15656 0 15716 88
use opamp  opamp_0 ~/tt06-fet-opamp/mag
timestamp 1713125316
transform -1 0 13182 0 -1 1498
box -1339 -2666 2810 300
<< labels >>
flabel metal4 s 15487 22476 15517 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 15855 22476 15885 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 15119 22476 15149 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15656 0 15716 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13448 0 13508 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11240 0 11300 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9032 0 9092 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 6824 0 6884 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 4616 0 4676 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 2408 0 2468 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 200 0 260 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 14751 22476 14781 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 14015 22476 14045 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13647 22476 13677 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12911 22476 12941 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12543 22476 12573 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11807 22476 11837 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11439 22476 11469 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10703 22476 10733 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10335 22476 10365 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9599 22476 9629 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9231 22476 9261 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 2975 22476 3005 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 2607 22476 2637 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 2239 22476 2269 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 1871 22476 1901 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 1503 22476 1533 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 1135 22476 1165 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 767 22476 797 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 399 22476 429 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 5919 22476 5949 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 5183 22476 5213 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 4815 22476 4845 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 4079 22476 4109 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 3711 22476 3741 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 8495 22476 8525 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8127 22476 8157 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 7391 22476 7421 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 7023 22476 7053 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 6287 22476 6317 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 250 22076 1 FreeSans 1 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 4900 1436 5050 22412 1 FreeSans 1 0 0 0 VGND
port 52 n
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
