magic
tech sky130A
magscale 1 2
timestamp 1713057736
<< nwell >>
rect -1199 -384 1199 384
<< pmos >>
rect -1003 -164 -803 236
rect -745 -164 -545 236
rect -487 -164 -287 236
rect -229 -164 -29 236
rect 29 -164 229 236
rect 287 -164 487 236
rect 545 -164 745 236
rect 803 -164 1003 236
<< pdiff >>
rect -1061 224 -1003 236
rect -1061 -152 -1049 224
rect -1015 -152 -1003 224
rect -1061 -164 -1003 -152
rect -803 224 -745 236
rect -803 -152 -791 224
rect -757 -152 -745 224
rect -803 -164 -745 -152
rect -545 224 -487 236
rect -545 -152 -533 224
rect -499 -152 -487 224
rect -545 -164 -487 -152
rect -287 224 -229 236
rect -287 -152 -275 224
rect -241 -152 -229 224
rect -287 -164 -229 -152
rect -29 224 29 236
rect -29 -152 -17 224
rect 17 -152 29 224
rect -29 -164 29 -152
rect 229 224 287 236
rect 229 -152 241 224
rect 275 -152 287 224
rect 229 -164 287 -152
rect 487 224 545 236
rect 487 -152 499 224
rect 533 -152 545 224
rect 487 -164 545 -152
rect 745 224 803 236
rect 745 -152 757 224
rect 791 -152 803 224
rect 745 -164 803 -152
rect 1003 224 1061 236
rect 1003 -152 1015 224
rect 1049 -152 1061 224
rect 1003 -164 1061 -152
<< pdiffc >>
rect -1049 -152 -1015 224
rect -791 -152 -757 224
rect -533 -152 -499 224
rect -275 -152 -241 224
rect -17 -152 17 224
rect 241 -152 275 224
rect 499 -152 533 224
rect 757 -152 791 224
rect 1015 -152 1049 224
<< nsubdiff >>
rect -1163 314 -1067 348
rect 1067 314 1163 348
rect -1163 -314 -1129 314
rect 1129 -314 1163 314
rect -1163 -348 1163 -314
<< nsubdiffcont >>
rect -1067 314 1067 348
<< poly >>
rect -1003 236 -803 262
rect -745 236 -545 262
rect -487 236 -287 262
rect -229 236 -29 262
rect 29 236 229 262
rect 287 236 487 262
rect 545 236 745 262
rect 803 236 1003 262
rect -1003 -211 -803 -164
rect -1003 -245 -987 -211
rect -819 -245 -803 -211
rect -1003 -261 -803 -245
rect -745 -211 -545 -164
rect -745 -245 -729 -211
rect -561 -245 -545 -211
rect -745 -261 -545 -245
rect -487 -211 -287 -164
rect -487 -245 -471 -211
rect -303 -245 -287 -211
rect -487 -261 -287 -245
rect -229 -211 -29 -164
rect -229 -245 -213 -211
rect -45 -245 -29 -211
rect -229 -261 -29 -245
rect 29 -211 229 -164
rect 29 -245 45 -211
rect 213 -245 229 -211
rect 29 -261 229 -245
rect 287 -211 487 -164
rect 287 -245 303 -211
rect 471 -245 487 -211
rect 287 -261 487 -245
rect 545 -211 745 -164
rect 545 -245 561 -211
rect 729 -245 745 -211
rect 545 -261 745 -245
rect 803 -211 1003 -164
rect 803 -245 819 -211
rect 987 -245 1003 -211
rect 803 -261 1003 -245
<< polycont >>
rect -987 -245 -819 -211
rect -729 -245 -561 -211
rect -471 -245 -303 -211
rect -213 -245 -45 -211
rect 45 -245 213 -211
rect 303 -245 471 -211
rect 561 -245 729 -211
rect 819 -245 987 -211
<< locali >>
rect -1163 -314 -1129 348
rect -1049 224 -1015 240
rect -1049 -168 -1015 -152
rect -791 224 -757 240
rect -791 -168 -757 -152
rect -533 224 -499 240
rect -533 -168 -499 -152
rect -275 224 -241 240
rect -275 -168 -241 -152
rect -17 224 17 240
rect -17 -168 17 -152
rect 241 224 275 240
rect 241 -168 275 -152
rect 499 224 533 240
rect 499 -168 533 -152
rect 757 224 791 240
rect 757 -168 791 -152
rect 1015 224 1049 240
rect 1015 -168 1049 -152
rect -1003 -245 -987 -211
rect -819 -245 -803 -211
rect -745 -245 -729 -211
rect -561 -245 -545 -211
rect -487 -245 -471 -211
rect -303 -245 -287 -211
rect -229 -245 -213 -211
rect -45 -245 -29 -211
rect 29 -245 45 -211
rect 213 -245 229 -211
rect 287 -245 303 -211
rect 471 -245 487 -211
rect 545 -245 561 -211
rect 729 -245 745 -211
rect 803 -245 819 -211
rect 987 -245 1003 -211
rect 1129 -314 1163 348
rect -1163 -348 1163 -314
<< viali >>
rect -1129 314 -1067 348
rect -1067 314 1067 348
rect 1067 314 1129 348
rect -1049 -152 -1015 224
rect -791 -152 -757 224
rect -533 -152 -499 224
rect -275 -152 -241 224
rect -17 -152 17 224
rect 241 -152 275 224
rect 499 -152 533 224
rect 757 -152 791 224
rect 1015 -152 1049 224
rect -987 -245 -819 -211
rect -729 -245 -561 -211
rect -471 -245 -303 -211
rect -213 -245 -45 -211
rect 45 -245 213 -211
rect 303 -245 471 -211
rect 561 -245 729 -211
rect 819 -245 987 -211
<< metal1 >>
rect -1141 348 1141 354
rect -1141 314 -1129 348
rect 1129 314 1141 348
rect -1141 308 1141 314
rect -1055 224 -1009 236
rect -1055 -152 -1049 224
rect -1015 -152 -1009 224
rect -1055 -164 -1009 -152
rect -797 224 -751 236
rect -797 -152 -791 224
rect -757 -152 -751 224
rect -797 -164 -751 -152
rect -539 224 -493 236
rect -539 -152 -533 224
rect -499 -152 -493 224
rect -539 -164 -493 -152
rect -281 224 -235 236
rect -281 -152 -275 224
rect -241 -152 -235 224
rect -281 -164 -235 -152
rect -23 224 23 236
rect -23 -152 -17 224
rect 17 -152 23 224
rect -23 -164 23 -152
rect 235 224 281 236
rect 235 -152 241 224
rect 275 -152 281 224
rect 235 -164 281 -152
rect 493 224 539 236
rect 493 -152 499 224
rect 533 -152 539 224
rect 493 -164 539 -152
rect 751 224 797 236
rect 751 -152 757 224
rect 791 -152 797 224
rect 751 -164 797 -152
rect 1009 224 1055 236
rect 1009 -152 1015 224
rect 1049 -152 1055 224
rect 1009 -164 1055 -152
rect -999 -211 -807 -205
rect -999 -245 -987 -211
rect -819 -245 -807 -211
rect -999 -251 -807 -245
rect -741 -211 -549 -205
rect -741 -245 -729 -211
rect -561 -245 -549 -211
rect -741 -251 -549 -245
rect -483 -211 -291 -205
rect -483 -245 -471 -211
rect -303 -245 -291 -211
rect -483 -251 -291 -245
rect -225 -211 -33 -205
rect -225 -245 -213 -211
rect -45 -245 -33 -211
rect -225 -251 -33 -245
rect 33 -211 225 -205
rect 33 -245 45 -211
rect 213 -245 225 -211
rect 33 -251 225 -245
rect 291 -211 483 -205
rect 291 -245 303 -211
rect 471 -245 483 -211
rect 291 -251 483 -245
rect 549 -211 741 -205
rect 549 -245 561 -211
rect 729 -245 741 -211
rect 549 -251 741 -245
rect 807 -211 999 -205
rect 807 -245 819 -211
rect 987 -245 999 -211
rect 807 -251 999 -245
<< properties >>
string FIXED_BBOX -1146 -331 1146 331
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
