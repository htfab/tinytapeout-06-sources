magic
tech sky130A
magscale 1 2
timestamp 1713540189
<< nwell >>
rect -425 -1819 425 1819
<< pmos >>
rect -229 -1600 -29 1600
rect 29 -1600 229 1600
<< pdiff >>
rect -287 1588 -229 1600
rect -287 -1588 -275 1588
rect -241 -1588 -229 1588
rect -287 -1600 -229 -1588
rect -29 1588 29 1600
rect -29 -1588 -17 1588
rect 17 -1588 29 1588
rect -29 -1600 29 -1588
rect 229 1588 287 1600
rect 229 -1588 241 1588
rect 275 -1588 287 1588
rect 229 -1600 287 -1588
<< pdiffc >>
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
<< nsubdiff >>
rect -389 1749 -293 1783
rect 293 1749 389 1783
rect -389 1687 -355 1749
rect 355 1687 389 1749
rect -389 -1749 -355 -1687
rect 355 -1749 389 -1687
rect -389 -1783 -293 -1749
rect 293 -1783 389 -1749
<< nsubdiffcont >>
rect -293 1749 293 1783
rect -389 -1687 -355 1687
rect 355 -1687 389 1687
rect -293 -1783 293 -1749
<< poly >>
rect -229 1681 -29 1697
rect -229 1647 -213 1681
rect -45 1647 -29 1681
rect -229 1600 -29 1647
rect 29 1681 229 1697
rect 29 1647 45 1681
rect 213 1647 229 1681
rect 29 1600 229 1647
rect -229 -1647 -29 -1600
rect -229 -1681 -213 -1647
rect -45 -1681 -29 -1647
rect -229 -1697 -29 -1681
rect 29 -1647 229 -1600
rect 29 -1681 45 -1647
rect 213 -1681 229 -1647
rect 29 -1697 229 -1681
<< polycont >>
rect -213 1647 -45 1681
rect 45 1647 213 1681
rect -213 -1681 -45 -1647
rect 45 -1681 213 -1647
<< locali >>
rect -389 1749 -293 1783
rect 293 1749 389 1783
rect -389 1687 -355 1749
rect 355 1687 389 1749
rect -229 1647 -213 1681
rect -45 1647 -29 1681
rect 29 1647 45 1681
rect 213 1647 229 1681
rect -275 1588 -241 1604
rect -275 -1604 -241 -1588
rect -17 1588 17 1604
rect -17 -1604 17 -1588
rect 241 1588 275 1604
rect 241 -1604 275 -1588
rect -229 -1681 -213 -1647
rect -45 -1681 -29 -1647
rect 29 -1681 45 -1647
rect 213 -1681 229 -1647
rect -389 -1749 -355 -1687
rect 355 -1749 389 -1687
rect -389 -1783 -293 -1749
rect 293 -1783 389 -1749
<< viali >>
rect -213 1647 -45 1681
rect 45 1647 213 1681
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
rect -213 -1681 -45 -1647
rect 45 -1681 213 -1647
<< metal1 >>
rect -225 1681 -33 1687
rect -225 1647 -213 1681
rect -45 1647 -33 1681
rect -225 1641 -33 1647
rect 33 1681 225 1687
rect 33 1647 45 1681
rect 213 1647 225 1681
rect 33 1641 225 1647
rect -281 1588 -235 1600
rect -281 -1588 -275 1588
rect -241 -1588 -235 1588
rect -281 -1600 -235 -1588
rect -23 1588 23 1600
rect -23 -1588 -17 1588
rect 17 -1588 23 1588
rect -23 -1600 23 -1588
rect 235 1588 281 1600
rect 235 -1588 241 1588
rect 275 -1588 281 1588
rect 235 -1600 281 -1588
rect -225 -1647 -33 -1641
rect -225 -1681 -213 -1647
rect -45 -1681 -33 -1647
rect -225 -1687 -33 -1681
rect 33 -1647 225 -1641
rect 33 -1681 45 -1647
rect 213 -1681 225 -1647
rect 33 -1687 225 -1681
<< properties >>
string FIXED_BBOX -372 -1766 372 1766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 16.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
