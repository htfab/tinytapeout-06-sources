magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< nwell >>
rect -1199 -419 1199 419
<< pmos >>
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
<< pdiff >>
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
<< pdiffc >>
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
<< nsubdiff >>
rect -1163 349 -1067 383
rect 1067 349 1163 383
rect -1163 -349 -1129 349
rect 1129 -349 1163 349
rect -1163 -383 1163 -349
<< nsubdiffcont >>
rect -1067 349 1067 383
<< poly >>
rect -1003 281 -803 297
rect -1003 247 -987 281
rect -819 247 -803 281
rect -1003 200 -803 247
rect -745 281 -545 297
rect -745 247 -729 281
rect -561 247 -545 281
rect -745 200 -545 247
rect -487 281 -287 297
rect -487 247 -471 281
rect -303 247 -287 281
rect -487 200 -287 247
rect -229 281 -29 297
rect -229 247 -213 281
rect -45 247 -29 281
rect -229 200 -29 247
rect 29 281 229 297
rect 29 247 45 281
rect 213 247 229 281
rect 29 200 229 247
rect 287 281 487 297
rect 287 247 303 281
rect 471 247 487 281
rect 287 200 487 247
rect 545 281 745 297
rect 545 247 561 281
rect 729 247 745 281
rect 545 200 745 247
rect 803 281 1003 297
rect 803 247 819 281
rect 987 247 1003 281
rect 803 200 1003 247
rect -1003 -247 -803 -200
rect -1003 -281 -987 -247
rect -819 -281 -803 -247
rect -1003 -297 -803 -281
rect -745 -247 -545 -200
rect -745 -281 -729 -247
rect -561 -281 -545 -247
rect -745 -297 -545 -281
rect -487 -247 -287 -200
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -487 -297 -287 -281
rect -229 -247 -29 -200
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect -229 -297 -29 -281
rect 29 -247 229 -200
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 29 -297 229 -281
rect 287 -247 487 -200
rect 287 -281 303 -247
rect 471 -281 487 -247
rect 287 -297 487 -281
rect 545 -247 745 -200
rect 545 -281 561 -247
rect 729 -281 745 -247
rect 545 -297 745 -281
rect 803 -247 1003 -200
rect 803 -281 819 -247
rect 987 -281 1003 -247
rect 803 -297 1003 -281
<< polycont >>
rect -987 247 -819 281
rect -729 247 -561 281
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect 561 247 729 281
rect 819 247 987 281
rect -987 -281 -819 -247
rect -729 -281 -561 -247
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
rect 561 -281 729 -247
rect 819 -281 987 -247
<< locali >>
rect -1163 -349 -1129 383
rect -1003 247 -987 281
rect -819 247 -803 281
rect -745 247 -729 281
rect -561 247 -545 281
rect -487 247 -471 281
rect -303 247 -287 281
rect -229 247 -213 281
rect -45 247 -29 281
rect 29 247 45 281
rect 213 247 229 281
rect 287 247 303 281
rect 471 247 487 281
rect 545 247 561 281
rect 729 247 745 281
rect 803 247 819 281
rect 987 247 1003 281
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect -1003 -281 -987 -247
rect -819 -281 -803 -247
rect -745 -281 -729 -247
rect -561 -281 -545 -247
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 287 -281 303 -247
rect 471 -281 487 -247
rect 545 -281 561 -247
rect 729 -281 745 -247
rect 803 -281 819 -247
rect 987 -281 1003 -247
rect 1129 -349 1163 383
rect -1163 -383 1163 -349
<< viali >>
rect -1129 349 -1067 383
rect -1067 349 1067 383
rect 1067 349 1129 383
rect -987 247 -819 281
rect -729 247 -561 281
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect 561 247 729 281
rect 819 247 987 281
rect -1049 -171 -1015 -21
rect -791 21 -757 171
rect -533 -171 -499 -21
rect -275 21 -241 171
rect -17 -171 17 -21
rect 241 21 275 171
rect 499 -171 533 -21
rect 757 21 791 171
rect 1015 -171 1049 -21
rect -987 -281 -819 -247
rect -729 -281 -561 -247
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
rect 561 -281 729 -247
rect 819 -281 987 -247
<< metal1 >>
rect -1141 383 1141 389
rect -1141 349 -1129 383
rect 1129 349 1141 383
rect -1141 343 1141 349
rect -999 281 -807 287
rect -999 247 -987 281
rect -819 247 -807 281
rect -999 241 -807 247
rect -741 281 -549 287
rect -741 247 -729 281
rect -561 247 -549 281
rect -741 241 -549 247
rect -483 281 -291 287
rect -483 247 -471 281
rect -303 247 -291 281
rect -483 241 -291 247
rect -225 281 -33 287
rect -225 247 -213 281
rect -45 247 -33 281
rect -225 241 -33 247
rect 33 281 225 287
rect 33 247 45 281
rect 213 247 225 281
rect 33 241 225 247
rect 291 281 483 287
rect 291 247 303 281
rect 471 247 483 281
rect 291 241 483 247
rect 549 281 741 287
rect 549 247 561 281
rect 729 247 741 281
rect 549 241 741 247
rect 807 281 999 287
rect 807 247 819 281
rect 987 247 999 281
rect 807 241 999 247
rect -797 171 -751 183
rect -797 21 -791 171
rect -757 21 -751 171
rect -797 9 -751 21
rect -281 171 -235 183
rect -281 21 -275 171
rect -241 21 -235 171
rect -281 9 -235 21
rect 235 171 281 183
rect 235 21 241 171
rect 275 21 281 171
rect 235 9 281 21
rect 751 171 797 183
rect 751 21 757 171
rect 791 21 797 171
rect 751 9 797 21
rect -1055 -21 -1009 -9
rect -1055 -171 -1049 -21
rect -1015 -171 -1009 -21
rect -1055 -183 -1009 -171
rect -539 -21 -493 -9
rect -539 -171 -533 -21
rect -499 -171 -493 -21
rect -539 -183 -493 -171
rect -23 -21 23 -9
rect -23 -171 -17 -21
rect 17 -171 23 -21
rect -23 -183 23 -171
rect 493 -21 539 -9
rect 493 -171 499 -21
rect 533 -171 539 -21
rect 493 -183 539 -171
rect 1009 -21 1055 -9
rect 1009 -171 1015 -21
rect 1049 -171 1055 -21
rect 1009 -183 1055 -171
rect -999 -247 -807 -241
rect -999 -281 -987 -247
rect -819 -281 -807 -247
rect -999 -287 -807 -281
rect -741 -247 -549 -241
rect -741 -281 -729 -247
rect -561 -281 -549 -247
rect -741 -287 -549 -281
rect -483 -247 -291 -241
rect -483 -281 -471 -247
rect -303 -281 -291 -247
rect -483 -287 -291 -281
rect -225 -247 -33 -241
rect -225 -281 -213 -247
rect -45 -281 -33 -247
rect -225 -287 -33 -281
rect 33 -247 225 -241
rect 33 -281 45 -247
rect 213 -281 225 -247
rect 33 -287 225 -281
rect 291 -247 483 -241
rect 291 -281 303 -247
rect 471 -281 483 -247
rect 291 -287 483 -281
rect 549 -247 741 -241
rect 549 -281 561 -247
rect 729 -281 741 -247
rect 549 -287 741 -281
rect 807 -247 999 -241
rect 807 -281 819 -247
rect 987 -281 999 -247
rect 807 -287 999 -281
<< properties >>
string FIXED_BBOX -1146 -366 1146 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
