* PEX produced on Sun Mar 10 05:48:33 PM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_hpretl_tt06_tempsens.ext - technology: sky130A

.subckt tt_um_hpretl_tt06_tempsens clk ena rst_n ui_in[2] ui_in[4] ui_in[6] uio_in[1]
+ uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[4] uio_oe[5] uio_oe[7]
+ uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[5] uo_out[6] uo_out[7] ui_in[1] uio_out[2] ui_in[3] uio_out[0] uio_oe[3]
+ uo_out[0] ui_in[5] uio_oe[1] uio_oe[6] ui_in[7] uio_oe[0] uio_out[1] uio_oe[2] uio_in[0]
+ ui_in[0] uo_out[4] uio_in[2] VPWR VGND
X0 a_5989_7669# a_5823_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=498 ps=4.72k w=0.87 l=4.73
X2 a_14935_1941# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_17051_1941# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_12531_9545# _107_ a_12449_9301# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 ts.ts_core.dac_vout_ana_ net14 a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 _051_ _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_17935_13363# net70 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 _099_ _098_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 VPWR net35 ts.ts_core.capload\[7\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR _062_ a_11679_6183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VPWR a_13327_9813# _089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND _070_ a_10686_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X15 a_11127_15797# a_10952_15823# a_11306_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X16 a_8653_3677# a_8175_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X17 VGND net7 a_13834_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND _154_ a_8625_4438# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X19 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=331 ps=3.4k w=0.55 l=4.73
X20 net19 a_8399_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 net14 a_17783_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_10969_6031# a_9779_6031# a_10860_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X23 ts.ts_core.dac_vout_ana_ net15 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_5081_4777# a_3891_4405# a_4972_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X25 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_3981_8449# a_3763_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X27 net69 a_18234_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 a_17051_1941# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X30 ts.ts_core.dac_vout_ana_ net14 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VPWR _112_ _114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VGND clknet_2_0__leaf_clk a_3247_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VGND net69 a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.dcdel_out_n VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X35 net9 a_18671_14451# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 _012_ _167_ a_1861_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X37 a_4588_5807# net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X38 VPWR a_17507_8751# a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X39 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X40 VGND net19 a_12489_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 VGND clknet_2_2__leaf_clk a_5823_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X42 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X43 VGND a_3854_3967# a_3812_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X44 a_4590_12381# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X45 a_12884_4777# a_11803_4405# a_12537_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X46 a_2869_10205# ts.ts_ctrl.temp_ctr\[7\] a_2787_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X47 a_14475_5205# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X49 a_13499_11247# a_13445_11159# a_13399_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X50 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X51 a_10335_4117# a_10147_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X52 a_17695_4399# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X53 a_14567_6575# a_14379_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X54 a_8856_10383# _055_ a_8468_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X55 VPWR a_16043_7271# a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X56 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X57 a_10023_4917# a_9848_4943# a_10202_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X58 a_1589_8725# a_1371_9129# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X59 a_17935_13363# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X60 a_9061_16665# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 VPWR _098_ a_13275_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X62 a_12851_7119# _111_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X63 ts.ts_core.dac_vout_ana_ net15 a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X64 a_9960_10383# ts.o_res\[8\] a_9770_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X65 _086_ a_8859_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X66 a_16569_1455# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X67 VPWR net9 a_8809_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X68 a_4111_4221# a_3413_3855# a_3854_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X69 VGND clknet_0_clk a_7838_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 VGND uio_out[2] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X70 _010_ _164_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 VGND net69 a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X72 a_8638_17821# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X73 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X74 a_6711_15657# a_6265_15285# a_6615_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X75 VPWR a_14663_5461# a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X76 VGND net53 a_1407_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X77 a_9850_4399# a_9577_4405# a_9765_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X78 _064_ a_13731_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X79 net10 a_18848_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X80 a_14475_6293# a_14287_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X81 a_12757_12015# _068_ a_12673_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X82 a_12819_2223# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X83 a_15591_5487# ts.ts_ctrl.state\[1\] _112_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X84 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X85 a_9464_16911# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X86 a_11969_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X87 a_12808_5603# ts.ts_ctrl.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.148 ps=1.34 w=0.42 l=0.15
X88 a_14195_9295# _135_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X89 a_2290_7119# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X90 a_8235_8790# ts.o_res\[3\] a_8235_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 VPWR clknet_2_3__leaf_clk a_11619_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X92 a_16687_9447# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X93 a_6945_11225# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X94 VGND a_4411_12319# a_4345_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X95 a_4503_4777# a_4057_4405# a_4407_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X96 VGND net9 a_8809_8534# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X97 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X98 a_11985_17429# a_11767_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X99 a_15304_8207# net47 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X100 a_9045_9839# ts.ts_ctrl.temp_ctr\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X101 a_16775_7663# a_16587_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X102 a_8657_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 a_3105_14557# a_3061_14165# a_2939_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X104 a_2695_12559# ts.ts_ctrl.temp_ctr\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X105 a_8749_12809# ts.o_res\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X106 VPWR a_9971_743# a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X107 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X109 a_12809_11247# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X110 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X112 a_6817_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X115 VGND net67 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X116 a_10689_12809# ts.o_res\[6\] a_10607_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X117 a_9333_17999# a_9298_18251# a_9095_17973# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X118 VGND net67 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X119 _135_ a_14177_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X120 a_7075_13481# a_6725_13109# a_6980_13469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X122 VGND net20 a_5773_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X123 a_7737_1455# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X124 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X125 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X126 a_10313_3855# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X127 a_16591_1135# a_16403_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X128 VGND _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X129 a_9687_10633# _075_ a_9770_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X130 VGND net67 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X131 net16 a_5423_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X133 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _065_ a_16170_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X134 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X135 VPWR net9 a_7521_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X136 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X137 a_4956_5461# _201_ a_5085_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X138 VPWR a_2111_11231# a_2098_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X140 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X141 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X142 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X143 ts.ts_core.dac_vout_ana_ net71 a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X144 a_6265_15285# a_6099_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X145 a_7321_16733# ts.ts_ctrl.temp_ctr\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X146 VGND a_11679_6183# _136_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X147 VPWR a_15399_12711# a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X148 ts.ts_core.dac_vout_ana_ net14 a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X149 a_10441_15577# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X150 _196_ ts.ts_ctrl.temp_ctr\[17\] a_3977_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X151 VPWR a_16955_4943# a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X152 VGND net68 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X153 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X154 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X155 a_3503_10927# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X156 a_4131_17833# a_3615_17461# a_4036_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X157 VPWR a_16127_591# a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X158 a_17695_6575# a_17507_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X159 VGND net9 a_7521_8534# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X160 a_1276_14735# _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X161 VPWR clknet_0_clk a_4986_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X163 VPWR a_16403_10383# a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X164 a_12997_6031# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X165 _059_ net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X166 VPWR ts.ts_ctrl.state\[0\] a_10605_3427# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X167 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X168 VPWR a_16687_9447# a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X169 uo_out[1] a_11456_11247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 a_8481_7119# ts.ts_ctrl.temp_ctr\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X171 VPWR a_9095_17973# ts.o_res\[12\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X172 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X173 a_10335_1941# a_10147_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X174 a_8179_5865# a_7663_5493# a_8084_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X175 a_16569_10383# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X176 ts.ts_core.dac_vout_ana_ net72 a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X177 net14 a_17783_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X178 net11 a_18756_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X179 VPWR net53 a_1407_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X180 VGND net67 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X181 VGND _112_ a_10227_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X182 _142_ a_18735_6059# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X183 _168_ a_2695_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X184 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X185 a_7759_1135# a_7571_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X186 VPWR _141_ a_18735_6059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
R1 uio_oe[0] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X188 a_17581_10159# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X189 uo_out[5] a_9524_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X190 VGND a_4495_16885# _018_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X192 a_10313_3855# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X193 VPWR a_9112_11989# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X194 VGND _083_ a_10585_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X195 a_4328_15823# a_3413_15823# a_3981_16065# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X196 a_13611_4917# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X197 a_17862_6281# _061_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X198 a_17121_4943# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X199 a_16591_10645# a_16403_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X200 VGND a_8632_16599# _214_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X201 a_13741_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13326_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X202 VPWR a_8459_17759# a_8446_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 VPWR a_7079_9055# a_7066_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X204 _019_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X205 a_1479_8751# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X206 a_18243_7983# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _096_ VGND sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X207 a_3517_12809# net62 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X208 a_1371_14735# a_855_14735# a_1276_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X209 VGND a_17332_3829# net67 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X210 VPWR clknet_2_0__leaf_clk net52 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X211 VPWR clknet_0_clk a_4513_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X212 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X214 a_9500_12015# _051_ a_9112_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X215 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X217 a_9353_12809# net8 a_9524_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R2 VGND uio_out[3] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X218 a_15212_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X219 a_6541_17999# a_6375_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X220 a_16477_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X221 VPWR _216_ a_10975_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X222 a_15741_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X223 a_8695_3553# clknet_2_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X224 VGND _184_ a_6457_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X225 a_7088_4777# a_6173_4405# a_6741_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X226 _119_ a_11343_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X227 a_14388_2223# a_15123_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X228 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X229 ts.ts_core.i_precharge_n a_13705_6353# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0986 ps=0.98 w=0.65 l=0.15
X230 a_12597_7663# _122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X231 a_14571_11623# net69 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X232 a_10401_4777# a_9411_4405# a_10275_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X233 a_15465_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X234 a_12507_17759# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X235 a_2131_14511# ts.ts_ctrl.temp_ctr\[9\] _175_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X236 VPWR ts.ts_ctrl.temp_ctr\[19\] _200_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X237 a_10068_13423# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X238 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X239 a_6461_591# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X240 a_3601_3855# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X241 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X242 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X243 a_15321_7663# _061_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X244 a_8491_7663# _090_ a_8573_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X245 a_11812_4105# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X246 a_9501_5185# a_9283_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X247 _059_ net11 a_14471_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 VGND a_4871_17759# ts.ts_ctrl.temp_ctr\[11\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X249 VGND net3 a_16354_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X250 VPWR a_4411_12319# a_4398_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X251 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X252 a_2755_8983# ts.ts_ctrl.temp_ctr\[2\] a_2929_9089# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X253 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X254 ts.ts_ctrl.temp_ctr\[15\] a_6251_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X255 a_9224_10927# _048_ a_8836_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X256 a_3663_15511# _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X257 VPWR a_6557_11713# a_6447_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X258 a_16960_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X259 a_4429_14557# ts.ts_ctrl.temp_ctr\[9\] a_4341_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X260 VGND net9 _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X261 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X262 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X263 a_10625_7352# ts.ts_ctrl.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X264 VPWR a_16311_12559# a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X265 a_5129_12559# a_5085_12801# a_4963_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X266 a_10011_3530# _202_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X267 VPWR _217_ a_9595_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X268 VGND net67 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X269 a_6839_853# a_6651_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X270 _061_ a_12047_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X272 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X274 a_8673_15253# a_8455_15657# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X275 VGND a_5893_17687# net63 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X276 VGND a_8447_6196# _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X277 _178_ _177_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X278 a_6631_9661# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X279 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X280 VPWR a_11803_1679# a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X281 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref _146_ a_18719_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X282 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X283 _112_ ts.ts_ctrl.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X284 VGND a_6607_17687# _183_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X285 a_4227_17833# a_3781_17461# a_4131_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X286 a_13869_3677# a_13825_3285# a_13703_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X287 a_14545_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X288 a_5140_15253# net58 a_5363_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X289 a_7075_13481# a_6559_13109# a_6980_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X290 VPWR clknet_2_1__leaf_clk net54 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X291 a_2290_11293# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X292 VPWR a_7640_13481# a_7815_13407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X293 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X294 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X295 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X296 a_12231_14735# a_11785_14735# a_12135_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X297 ts.ts_ctrl.temp_ctr\[18\] a_4687_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X298 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X299 VGND _047_ a_9716_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X300 a_9236_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X301 _038_ a_8767_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X303 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X304 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X305 a_17673_15599# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X306 a_10141_6575# ts.ts_ctrl.temp_ctr\[1\] _158_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X307 VPWR clknet_2_0__leaf_clk a_3891_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X308 a_15451_14423# net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X309 VPWR net9 a_12752_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X310 VGND _143_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X311 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
R3 ts.ts_core.capload\[2\].cap_30.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X312 a_2111_9055# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X313 _143_ _122_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X314 VGND a_11272_11471# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X315 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X316 a_6792_7271# ts.ts_ctrl.temp_ctr\[2\] a_6934_7446# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X317 a_12227_15657# a_11877_15285# a_12132_15645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X318 a_15948_9295# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X319 a_8941_13103# _085_ a_8859_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X320 VPWR _066_ a_10055_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X321 VGND _075_ a_8193_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X322 VPWR a_18335_2223# net72 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X323 VPWR a_14937_9955# _095_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.5 as=0.135 ps=1.27 w=1 l=0.15
X324 a_9643_14410# _208_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X325 VPWR a_17507_15279# a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X326 VGND a_18234_10927# net69 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 VPWR a_9800_13423# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 a_9629_13103# ts.o_res\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X329 a_14107_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X330 VGND net67 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X331 VPWR a_6904_8041# a_7079_7967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X332 a_10516_10633# ts.o_res\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X333 ts.o_res\[17\] a_7263_6879# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X334 _125_ a_12079_8457# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X335 VPWR a_13546_13335# _082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X336 a_11875_17455# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X337 a_8496_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X338 a_11847_16911# ts.ts_ctrl.temp_ctr\[13\] a_11484_17063# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X339 VGND a_2111_11231# a_2045_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X340 a_3413_10633# _170_ a_3329_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X341 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X342 a_12797_2543# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X343 a_9848_4943# a_8933_4943# a_9501_5185# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X344 a_15399_12711# net70 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X345 a_14471_8207# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X346 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X347 a_6435_11471# a_5989_11471# a_6339_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X348 VPWR a_9227_1135# a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X349 VPWR a_6515_6196# _044_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X350 _126_ a_10147_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X351 a_16315_5487# a_16127_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X352 a_17143_14191# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X353 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X354 a_7737_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X355 a_16315_853# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X356 a_8816_6183# ts.o_res\[1\] a_8958_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X357 VGND net68 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X358 net67 a_17332_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X359 a_16131_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X360 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X361 a_7252_12711# ts.o_res\[5\] a_7394_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X362 net65 a_15571_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X363 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X364 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X365 a_2305_10535# a_2401_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X366 a_6553_1455# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X367 a_13560_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X368 a_2859_5487# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X369 _202_ a_8879_4438# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X370 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X371 a_14388_2223# a_15123_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X372 a_7263_9269# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X373 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X374 a_9339_18582# ts.ts_ctrl.temp_ctr\[12\] a_9339_18909# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X375 VGND net67 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X376 a_9393_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X377 VGND net18 a_3105_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X378 a_10200_6031# _008_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X379 a_8105_15285# a_7939_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X380 VGND net67 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X381 VPWR _062_ _110_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X382 _069_ _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X383 VGND ts.ts_ctrl.temp_ctr\[10\] a_3944_14709# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X384 a_10233_16911# a_9043_16911# a_10124_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X385 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _061_ a_15321_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X386 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10147_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X387 a_16354_9071# _065_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X388 ts.ts_core.dac_vout_ana_ net47 a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 VGND net19 a_12029_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X390 a_4674_5309# a_3597_4943# a_4512_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X391 a_9556_14735# _033_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X392 a_12797_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X393 a_14384_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X394 a_12819_2223# a_12631_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X395 a_1501_8457# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X396 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X397 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X398 net9 a_18671_14451# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X399 VGND ts.ts_core.dcdel_capnode_ana_ a_11793_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X400 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X401 a_12875_14709# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X402 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X403 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X404 a_1276_12559# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X405 a_17143_7381# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X406 VGND a_7313_6005# a_7247_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X407 net70 a_17935_13363# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X408 a_6244_8029# _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X409 a_4490_8573# a_3413_8207# a_4328_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X410 a_3061_14165# a_2843_14569# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X411 _188_ _177_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X412 VPWR _094_ a_18325_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X413 ts.ts_core.dac_vout_ana_ net14 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X414 a_8657_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X415 VGND _067_ _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
R4 ts.ts_core.dac.vdac_single.einvp_batch\[0\].vref_38.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X417 ts.o_res\[13\] a_12507_17759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X418 a_10011_3530# _202_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X419 _091_ a_9770_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X420 _006_ a_16298_4719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X421 VPWR a_3316_5865# a_3491_5791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X422 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X423 a_7393_16733# ts.ts_ctrl.temp_ctr\[12\] a_7321_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X424 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X425 a_10335_3029# a_10147_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X426 a_15212_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X427 a_7381_1455# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X428 _200_ ts.ts_ctrl.temp_ctr\[19\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X429 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X430 a_16591_10645# a_16403_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X431 a_16315_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X432 a_9232_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X434 a_8468_10357# net8 a_8856_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X435 VPWR a_9235_1831# a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X436 VGND a_14717_9545# uio_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X437 VGND clknet_2_1__leaf_clk a_6007_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X438 VPWR ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_17783_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X439 a_4702_6031# ts.ts_ctrl.temp_ctr\[18\] a_4617_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X440 a_11797_6895# _109_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X441 a_10984_2223# a_11719_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X442 ts.ts_core.dac_vout_ana_ net14 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X443 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X444 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X445 a_2111_9055# a_1936_9129# a_2290_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X446 a_9651_14735# a_9135_14735# a_9556_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X447 a_15741_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X448 a_16683_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X449 VGND a_12157_13799# _056_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X451 VPWR _071_ a_10689_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X452 a_4871_17759# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X453 a_4952_11159# ts.o_res\[4\] a_5094_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X454 _049_ a_8386_11247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X455 VGND a_14584_8751# uio_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X456 ts.ts_core.dac_vout_ana_ net15 a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X457 a_13832_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X458 a_13556_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X459 VPWR a_12079_1135# a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X460 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X461 a_11969_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X462 a_9393_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X463 a_11969_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 a_6891_17999# a_6541_17999# a_6796_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X465 VGND _217_ a_9595_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X466 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X467 ts.ts_core.dac_vout_ana_ net14 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X468 a_8399_7369# _090_ a_8481_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X469 a_8448_9447# ts.o_res\[16\] a_8590_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X470 VPWR a_11760_14423# _212_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X471 ts.ts_core.capload\[2\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X472 ts.ts_core.dac_vout_ana_ net71 a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X473 VPWR a_14857_14342# a_14526_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X474 VPWR ts.ts_ctrl.temp_ctr\[4\] a_2695_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X475 a_13705_6353# a_13769_6296# a_13551_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X476 a_12353_14977# a_12135_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X477 a_9393_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X478 VPWR net3 a_16793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X479 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X480 a_16354_9071# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X481 VPWR a_11127_15797# a_11114_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X482 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X483 VGND ts.o_res\[13\] a_12157_13799# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X484 ts.ts_core.dac_vout_ana_ net72 a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X485 a_2397_15511# a_2493_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X487 VGND a_12127_7093# uio_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 _030_ a_5363_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X489 net4 a_18278_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X490 a_11119_4373# a_11478_4373# a_11255_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X491 ts.ts_core.dac_vout_ana_ net72 a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X493 a_11808_3855# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X494 VGND _137_ _190_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X495 a_17143_8469# a_16955_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X496 _020_ a_6690_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X497 a_12224_4765# _005_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X498 VPWR clknet_0_clk a_8022_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X499 VGND _077_ a_12896_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X500 _038_ a_8767_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X501 VPWR a_7815_4917# _211_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X502 a_6839_853# a_6651_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X503 VGND a_8695_3553# a_8656_3427# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X504 VPWR a_16043_8359# a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X505 a_2656_5853# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X506 a_11812_5193# a_12547_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X507 a_12946_13103# ts.o_res\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X508 VPWR a_10299_16885# a_10286_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 a_1585_10383# net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X510 a_18937_7147# _148_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X511 a_2098_10927# a_1021_10933# a_1936_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X512 a_17673_9071# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X513 a_11236_9295# _109_ a_10975_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X514 a_8360_15645# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X515 VPWR a_5179_16367# _138_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X516 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X517 VGND a_10299_16885# a_10233_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X518 a_8194_2223# a_7921_2229# a_8109_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X519 a_9415_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X520 VGND a_18671_14451# net9 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X521 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X522 ts.ts_core.capload\[13\].cap.Y net26 a_6185_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X523 a_2045_11305# a_855_10933# a_1936_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X524 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X525 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X526 VPWR a_4956_5461# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X527 VPWR a_2111_9055# a_2098_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X528 VPWR a_5515_10357# a_5502_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X529 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 VGND _074_ a_13503_10145# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X531 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X532 VGND net16 a_3013_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X533 VPWR _069_ a_12679_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X534 a_14913_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X535 VPWR _051_ a_11285_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X536 VPWR clknet_2_1__leaf_clk a_7663_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X537 VGND _193_ _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X538 a_6557_11713# a_6339_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X539 VPWR a_11803_2767# a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X540 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X541 _114_ _112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X542 VPWR a_6209_8181# a_6239_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X543 a_1021_10933# a_855_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X544 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X545 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X546 VPWR a_12056_3689# a_12231_3615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X547 VPWR a_14172_3689# a_14347_3615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X548 a_13553_12381# _073_ a_13453_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X549 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X550 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X551 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X552 VPWR _168_ a_2787_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X553 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X554 VGND ts.o_res\[14\] a_10961_13799# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X555 VPWR a_8491_2767# a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X557 VGND a_7815_4917# _211_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X558 VPWR a_11456_11247# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X559 VPWR a_7067_13812# _032_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X560 a_9415_2223# a_9227_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X561 ts.o_res\[15\] a_9195_15583# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X562 a_3413_3311# a_3177_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X564 a_3583_14495# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X565 VGND a_9643_14410# _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X566 a_7067_13812# _207_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X567 VGND a_8836_10901# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X568 VGND _131_ a_8583_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X569 ts.ts_core.dac_vout_ana_ net14 a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X570 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X571 a_13555_10901# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X572 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X573 a_10605_10383# _071_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X574 a_11285_10927# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X575 VPWR a_14287_4943# a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X576 a_1858_8207# _159_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X577 VGND a_9524_12559# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X578 a_9524_12559# ts.o_res\[5\] a_9440_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 VGND clknet_2_3__leaf_clk a_7203_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X580 a_7711_12886# ts.o_res\[5\] a_7252_12711# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X581 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X582 VPWR a_3981_8449# a_3871_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X583 VGND net70 a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X584 a_4772_12559# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X585 a_10335_3029# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X586 a_8500_1929# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X587 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X588 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X589 a_8446_17455# a_7369_17461# a_8284_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X590 a_15465_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X591 VGND _049_ a_9306_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X592 ts.ts_core.dac_vout_ana_ net14 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X593 a_17143_14191# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X594 a_3597_4943# a_3431_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X595 VPWR a_17507_8751# a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X596 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X597 a_7061_3855# a_7017_4097# a_6895_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X598 VGND a_7681_12533# a_7615_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X599 VPWR net61 a_1854_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X600 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X601 uio_out[5] a_14584_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X602 VPWR a_7263_9269# a_7250_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X603 a_3960_11305# a_2879_10933# a_3613_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X604 a_4312_4765# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X605 VPWR _189_ a_5269_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X606 VPWR net17 a_8996_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X607 a_15031_4373# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X608 VPWR clknet_2_3__leaf_clk a_6375_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X609 a_14475_5205# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X610 a_17143_7381# a_16955_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X611 a_3668_8207# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X612 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X613 a_6457_16911# _177_ _185_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X614 a_18847_14709# uio_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X615 a_15487_13909# a_15299_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X616 VGND a_6983_15797# a_6725_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X617 VPWR _047_ a_9500_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X618 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X619 VPWR a_16043_7271# a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X620 a_4057_4405# a_3891_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X621 a_6173_4405# a_6007_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X622 a_6880_16911# _185_ a_6780_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.114 ps=1 w=0.65 l=0.15
X623 a_12851_7119# _125_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X624 a_17877_9545# net3 a_17753_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.235 ps=1.47 w=1 l=0.15
X625 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 a_10980_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X627 VGND _211_ a_9560_18909# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X628 a_11396_3677# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X629 a_13512_3677# _006_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X630 ts.ts_core.dac_vout_ana_ net15 a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X631 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X632 a_16569_1455# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 VGND _066_ a_14453_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X634 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X636 a_6244_8029# _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X637 a_4398_12015# a_3321_12021# a_4236_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X639 ts.ts_ctrl.temp_ctr\[11\] a_4871_17759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X640 a_8657_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X641 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X642 a_8836_10901# _049_ a_9224_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X643 a_12819_2223# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X644 a_9236_841# a_9971_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X645 a_15259_13423# net12 a_14901_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X646 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X647 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X648 VPWR a_7456_17999# a_7631_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X649 a_12679_10071# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.34 w=0.42 l=0.15
X650 _047_ net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X651 VGND net67 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X652 ts.ts_ctrl.temp_ctr\[19\] a_5147_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X653 VPWR a_16495_10927# a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X654 VPWR a_15299_13647# a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X655 VGND net70 a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X656 VPWR a_15951_2919# a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X657 a_14085_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X658 a_9214_10159# _129_ a_9045_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X659 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_18755_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X660 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X661 a_16775_7663# a_16587_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X662 a_3977_6895# _194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X664 a_11975_5461# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X665 a_7815_4917# _153_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X666 ts.ts_ctrl.temp_ctr\[5\] a_2111_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X667 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X668 VGND _059_ _122_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X669 a_13959_13423# a_13905_13335# a_13859_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X670 _039_ a_9871_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X671 VGND net67 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X672 a_10294_7093# a_10147_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.331 ps=1.71 w=0.42 l=0.15
X673 VGND a_6516_11159# _209_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X674 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X675 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X676 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X677 a_11853_6059# _112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X679 VGND a_4329_13335# net62 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X680 ts.ts_core.dac_vout_ana_ net14 a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X681 a_4122_10927# a_3045_10933# a_3960_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X682 VGND net67 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X683 a_16960_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X684 a_15952_9545# a_16687_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X685 a_17673_15599# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X686 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X687 a_7737_1455# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X688 VGND net65 a_16298_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X689 a_2939_14569# a_2493_14197# a_2843_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X690 a_16964_13897# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X691 a_14296_4399# a_15031_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X692 VPWR net70 a_15299_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X693 a_5893_17687# a_5989_17429# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X694 a_9224_10927# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X695 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X696 a_14843_13621# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
R5 uio_oe[7] VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X697 VGND net68 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X698 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X699 VPWR a_14663_5461# a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X700 a_11863_17833# a_11417_17461# a_11767_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X701 a_11119_4373# ts.ts_ctrl.state\[1\] a_11338_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X702 ts.ts_core.capload\[5\].cap.Y net33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X703 a_11467_5825# _146_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X704 a_14475_6293# a_14287_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X705 a_12403_10177# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X706 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X708 ts.ts_core.dac_vout_ana_ net71 a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X709 VGND a_5381_11225# a_5315_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X710 a_14195_9295# _097_ a_14717_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X711 VGND a_18234_10927# net69 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X712 a_6430_14735# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X714 VGND _162_ a_2537_9323# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X715 a_11709_3285# a_11491_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X716 VPWR a_16955_4943# a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X718 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X719 VGND net68 a_14287_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X720 VPWR _151_ a_13551_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R6 VPWR tt_um_hpretl_tt06_tempsens_39.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X721 VPWR a_5423_4917# net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X722 a_16170_6895# _065_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X723 a_13399_11247# _068_ a_13295_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X724 VGND net68 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X725 ts.ts_core.dac_vout_ana_ net15 a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X726 a_6447_11837# a_5823_11471# a_6339_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X727 VPWR a_8362_2197# a_8289_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X728 a_4111_4221# a_3247_3855# a_3854_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X729 uo_out[6] a_9800_13423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X730 VPWR _047_ a_9629_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X731 VPWR a_13059_4703# ts.ts_ctrl.state\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X732 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X733 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X734 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X736 a_6523_4777# a_6173_4405# a_6428_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X737 a_7159_16599# ts.ts_ctrl.temp_ctr\[11\] a_7393_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X738 a_3583_14495# a_3408_14569# a_3762_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X739 a_6067_14191# _187_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X740 VGND clknet_2_3__leaf_clk a_7939_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X742 a_3329_10633# _172_ _014_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X743 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X744 a_14015_13077# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X746 VPWR a_9460_13799# _208_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X747 a_1775_8457# ts.ts_ctrl.temp_ctr\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X748 VPWR net11 a_13967_12711# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X749 VPWR a_4126_8983# _194_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X750 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X751 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X752 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X753 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X754 a_14935_1941# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X755 VGND ui_in[2] a_18278_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X756 a_17051_1941# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X757 VPWR _194_ a_4075_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X758 VGND a_3307_13799# _173_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X759 VPWR a_7088_6953# a_7263_6879# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X760 VGND a_6247_5461# a_5989_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X761 a_16293_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X762 a_5989_8757# a_5823_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X763 a_7088_9295# a_6173_9295# a_6741_9537# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X764 ts.ts_core.dac_vout_ana_ net15 a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X765 VPWR a_1589_12801# a_1479_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X766 VPWR a_10860_6031# a_11035_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X767 _067_ a_16180_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X768 a_17121_4943# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X769 a_7815_13407# a_7640_13481# a_7994_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X770 a_10138_11247# ts.o_res\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X771 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X772 VPWR a_18836_12711# a_18787_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.183 ps=1.37 w=1 l=0.15
X773 a_10335_4117# a_10147_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X774 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X775 a_18243_7983# _095_ _096_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X776 a_17695_4399# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X777 ts.ts_core.dac_vout_ana_ net14 a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R7 VGND net26 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X778 a_17695_6575# a_17507_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X779 VPWR net5 a_17862_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X780 a_15741_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X781 ts.ts_core.dac_vout_ana_ net14 a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X782 ts.ts_core.dac_vout_ana_ net71 a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X783 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X784 VPWR a_4683_13077# a_4425_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X785 a_17695_4399# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X786 a_14567_6575# a_14379_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X787 a_17599_6031# _065_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X788 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X789 a_9379_4943# a_8933_4943# a_9283_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X790 a_8532_11721# ts.o_res\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X791 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X792 VPWR _059_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X793 a_16771_10159# _065_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R8 net29 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X794 a_12056_3689# a_10975_3317# a_11709_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X795 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X796 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X797 VPWR a_15943_6031# a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X798 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X799 a_17862_6281# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X800 a_15304_8207# net47 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X801 VPWR a_6651_591# a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X802 a_14526_14165# a_14379_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.331 ps=1.71 w=0.42 l=0.15
X803 _069_ _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X804 VGND _216_ a_10975_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X805 _198_ a_4075_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X806 VPWR _114_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X807 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X808 a_6631_4399# a_6007_4405# a_6523_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X809 a_8155_4737# _139_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X810 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X811 VGND _115_ a_12079_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X812 a_15948_9295# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X813 a_16661_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X814 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X815 VPWR net55 a_9411_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X816 VGND a_8399_18543# net8 VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X817 VPWR ts.ts_ctrl.temp_ctr\[9\] a_4259_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X818 VGND clknet_2_0__leaf_clk a_855_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X819 VPWR ts.ts_ctrl.temp_ctr\[0\] a_10141_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X820 _048_ a_8532_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X821 _138_ a_5179_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X822 VPWR net6 a_15321_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X823 VGND a_13967_12711# _088_ VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X824 a_10313_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X825 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X826 a_2609_12381# ts.ts_ctrl.temp_ctr\[5\] a_2537_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X827 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
R9 VPWR tt_um_hpretl_tt06_tempsens_42.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X828 a_8856_10383# _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X829 VPWR a_10391_14709# a_10378_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X830 VPWR a_2305_10535# net60 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X831 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X833 a_18821_6059# _139_ a_18735_6059# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X834 VGND _075_ a_8837_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X835 VPWR a_16495_12015# a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X836 VGND a_12047_6835# _061_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X837 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X838 a_12853_12015# _073_ a_12757_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X839 _163_ a_2451_9323# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X840 VGND a_12967_15583# a_12901_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X841 VPWR _059_ _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X843 ts.ts_core.capload\[3\].cap.Y net31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X844 VPWR net67 a_7571_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X845 a_10585_13647# ts.ts_ctrl.temp_ctr\[6\] a_10239_13897# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X846 a_6998_17161# _183_ a_6690_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.22 ps=1.44 w=1 l=0.15
X847 VGND net52 a_3247_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X848 a_9415_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X849 a_16569_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X850 VGND a_8362_2197# a_8320_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X851 VPWR a_7681_12533# a_7711_12886# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X852 _075_ a_14707_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X853 _139_ a_12597_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.172 ps=1.35 w=1 l=0.15
X854 a_13183_7983# _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X855 a_3641_6941# _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X856 VGND a_3299_9269# _164_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X857 VGND a_8851_3285# a_8782_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X858 a_3763_8207# a_3247_8207# a_3668_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X859 a_12123_14557# ts.ts_ctrl.temp_ctr\[9\] a_11760_14423# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X860 a_17051_14997# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X862 a_11059_9955# _092_ a_10977_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X863 a_15948_9295# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X864 a_9235_1831# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X865 VPWR a_15299_13647# a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X866 a_6615_15657# a_6265_15285# a_6520_15645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X867 a_6428_6941# _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X868 VPWR clknet_2_0__leaf_clk a_6007_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X869 a_5607_12533# a_5432_12559# a_5786_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X870 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd a_18335_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X871 uio_out[7] a_14717_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X872 a_1762_14191# _173_ a_1459_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X873 a_14107_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X874 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X875 a_16465_5193# _098_ a_16393_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X876 _127_ a_10138_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X877 VGND a_11035_6005# a_10969_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X878 VPWR a_12231_3615# ts.ts_ctrl.state\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X879 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X880 a_1775_12015# ts.ts_ctrl.temp_ctr\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X881 VPWR a_11803_1679# a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X882 a_10313_3855# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X883 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X884 a_10286_17277# a_9209_16911# a_10124_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X885 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X886 a_1585_11721# _164_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X887 VGND _164_ a_1585_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X888 VGND a_18671_14451# net9 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X889 VGND a_12157_9813# _070_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X890 a_6238_15101# a_5161_14735# a_6076_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X891 a_12267_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X892 VPWR a_9227_1135# a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X893 VPWR a_18753_10548# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X895 a_16315_853# a_16127_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X896 ts.ts_core.capload\[8\].cap.Y net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X897 VPWR a_15575_3855# a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X898 a_16315_5487# a_16127_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X899 a_6741_6549# a_6523_6953# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X900 ts.ts_core.dac_vout_ana_ net72 a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X901 ts.ts_core.dac_vout_ana_ net15 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X902 VGND net68 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X903 a_6629_15975# a_6725_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X904 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X905 ts.ts_ctrl.state\[1\] a_13059_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X906 a_6987_17999# a_6541_17999# a_6891_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X907 VPWR a_9771_18236# a_9702_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X908 a_7759_1135# a_7571_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X909 a_16683_10927# a_16495_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X911 a_10313_3855# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X912 a_11597_13423# ts.ts_ctrl.temp_ctr\[10\] a_11159_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X913 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X914 VGND a_6515_6196# _044_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X915 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X916 a_18293_4020# ui_in[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X917 a_13101_7369# _125_ a_12127_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X918 _135_ a_14177_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X919 ts.o_res\[6\] a_10391_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X920 a_16293_13423# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X922 a_13551_8751# ts.ts_ctrl.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X923 a_17581_10159# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X924 a_15187_9955# _073_ a_15115_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X925 VGND a_11053_5719# _153_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X926 a_14935_1941# a_14747_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X927 a_17051_1941# a_16863_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X928 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X929 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X930 VGND a_17332_3829# net67 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X931 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X932 a_14388_2223# a_15123_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X933 VPWR a_6515_10058# _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X934 VGND _074_ a_14857_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X935 a_1633_14735# a_1589_14977# a_1467_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X936 VGND net67 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X937 a_10334_18365# a_9576_18267# a_9771_18236# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X938 _140_ net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.176 ps=1.39 w=1 l=0.15
X939 a_11808_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X940 a_5340_10383# a_4425_10383# a_4993_10625# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X941 ts.ts_ctrl.state\[0\] a_12231_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X942 ts.ts_ctrl.state\[2\] a_14347_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X943 VPWR a_4680_11445# net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X944 VGND a_11399_1109# a_11141_1109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X945 a_17783_5487# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 VGND a_9340_11471# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X947 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X948 a_11022_6397# a_9945_6031# a_10860_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X949 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X950 VPWR net52 a_3247_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X951 a_11812_4105# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X952 a_7159_16599# ts.ts_ctrl.temp_ctr\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X953 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X955 a_7387_17161# ts.ts_ctrl.temp_ctr\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X956 a_16293_591# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X957 VGND a_3479_6807# _197_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X958 VGND a_18774_3311# a_18880_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X959 a_4986_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X960 a_12946_13103# ts.o_res\[13\] a_12789_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X961 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X962 a_12901_15657# a_11711_15285# a_12792_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X963 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X964 VGND net69 a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X966 a_7624_17821# _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X967 a_7989_8534# ts.o_res\[2\] a_7775_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X968 a_11456_11247# _052_ a_11285_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X969 VGND a_8836_10901# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X970 VGND net70 a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X971 a_9792_12559# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X972 a_17143_7381# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X973 a_14857_10383# _073_ a_15125_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X974 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X975 a_12228_15823# ts.o_res\[10\] a_12007_16150# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X976 a_8590_3855# _153_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X977 a_15321_7663# _061_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X978 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X979 a_4513_13621# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X980 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X981 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _065_ a_16354_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X983 a_10984_2223# a_11719_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
R10 ts.ts_core.dac.vdac_single.einvp_batch\[0\].pupd_47.LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X984 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X985 VPWR ts.ts_ctrl.temp_ctr\[12\] a_7159_16599# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X986 a_13928_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X987 a_5167_16911# ts.ts_ctrl.temp_ctr\[11\] _181_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X988 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X989 a_7929_12335# ts.ts_ctrl.temp_ctr\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X990 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X991 a_15315_10383# a_15535_10357# _094_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X992 a_15212_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X993 VPWR a_15299_13647# a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X994 _061_ a_12047_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X995 a_12631_8457# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X996 a_7539_3829# a_7364_3855# a_7718_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X997 VGND net69 a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X998 VPWR a_2111_14709# ts.ts_ctrl.temp_ctr\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X999 VPWR clknet_2_0__leaf_clk a_2235_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1001 a_11478_4373# _110_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1002 a_7088_6953# a_6007_6581# a_6741_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1003 a_10607_12809# _088_ a_10689_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1004 a_10984_2223# a_11719_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1005 VGND ts.ts_ctrl.state\[0\] a_10147_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1006 _085_ a_7847_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1007 a_18234_10927# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1008 a_8851_3285# a_8656_3427# a_9161_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X1009 a_17143_14191# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1010 VGND a_5232_6005# _199_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X1011 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_15483_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1012 VGND net70 a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1013 a_15741_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1014 a_10570_14735# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1015 a_13183_7983# _113_ a_13601_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1016 VPWR a_18243_1135# net71 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R11 VGND net34 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1017 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1018 VGND a_14584_8751# uio_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1019 VPWR a_12079_1135# a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1020 a_11969_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1021 a_13921_6941# _113_ a_13821_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1022 _030_ a_5363_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1023 a_5780_8359# ts.ts_ctrl.temp_ctr\[3\] a_5922_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1024 a_16683_10927# a_16495_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1025 a_8179_5865# a_7829_5493# a_8084_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1027 a_9765_4399# net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1028 ts.ts_core.dcdel_capnode_ana_ ts.ts_core.i_precharge_n a_13892_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.183 ps=1.37 w=1 l=0.15
X1029 a_17695_8751# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1030 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1031 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1032 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1033 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1034 a_8399_7369# _090_ a_8481_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1035 a_3668_15823# _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
R12 VPWR tt_um_hpretl_tt06_tempsens_40.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1036 a_7640_13481# a_6559_13109# a_7293_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1037 VGND a_14063_10901# _077_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1038 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1039 a_8448_15975# ts.o_res\[15\] a_8590_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1040 a_16187_7895# _059_ a_16361_8001# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1042 VPWR a_6651_591# a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1044 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1045 ts.ts_core.dac_vout_ana_ net14 a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X1046 a_6427_16341# _114_ a_6858_16687# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X1047 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1048 _137_ a_6059_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1049 VGND _190_ a_5140_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X1050 a_14471_8207# _059_ _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1051 a_7171_13481# a_6725_13109# a_7075_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1052 VGND _173_ a_2131_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1053 a_7369_17461# a_7203_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1054 VPWR a_7180_15657# a_7355_15583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1055 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1056 VGND net69 a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1057 a_11808_3855# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1058 a_11057_9117# ts.ts_ctrl.state\[2\] a_10975_8864# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1059 VGND net70 a_17507_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1060 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14747_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1061 a_17143_8469# a_16955_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1062 a_8109_2223# ts.ts_core.tempdelay_async VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1063 ts.ts_core.dac_vout_ana_ net15 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1064 a_15671_11733# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1065 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1066 VGND _061_ a_16354_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1068 VPWR ts.o_res\[0\] a_9224_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1069 _117_ a_10607_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1070 _211_ a_7815_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1071 VGND a_5871_13335# _192_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1073 _053_ a_7775_8534# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1074 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref a_18234_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1075 net71 a_18243_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1076 _143_ _122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X1077 a_14567_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1078 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1079 ts.ts_core.dac_vout_ana_ net15 a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1080 a_4490_16189# a_3413_15823# a_4328_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1082 VGND a_4687_4917# a_4621_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1083 VGND a_7719_15797# a_7461_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X1084 a_8022_6575# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1085 VGND clk a_7286_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1086 VPWR a_7313_6005# a_7343_6358# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1087 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1088 a_4329_13335# a_4425_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X1089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1090 a_10023_4917# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1091 VPWR a_16955_14191# a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
R13 ts.ts_core.capload\[7\].cap_35.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1092 VGND net69 a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1093 a_11306_15823# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1094 a_2111_14709# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1095 VPWR net37 ts.ts_core.capload\[9\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1096 a_6921_2767# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1097 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1098 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1099 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1100 VGND a_15943_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1101 ts.ts_core.dac_vout_ana_ net14 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1102 a_8362_2197# a_8194_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1103 a_6067_14191# _189_ a_5975_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X1104 a_11437_7369# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1105 VPWR a_8284_17833# a_8459_17759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1106 a_12410_3677# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1107 a_4209_4943# a_4165_5185# a_4043_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1108 VPWR a_5780_8359# _205_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1109 a_5361_6031# _194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X1110 VPWR a_2659_10357# a_2401_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X1111 a_5922_8534# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1113 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1114 VGND a_11913_16885# a_11847_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1115 a_13892_1929# a_13643_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.321 ps=1.68 w=1 l=0.15
X1116 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1117 VGND a_7263_4703# a_7197_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1118 VGND a_5147_4703# a_5081_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1119 a_7066_7663# a_5989_7669# a_6904_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1120 ts.ts_core.dac_vout_ana_ net47 a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1121 a_11272_11471# _053_ a_11540_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1122 a_14717_9545# _097_ a_14195_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X1123 a_2271_4221# a_1573_3855# a_2014_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1124 a_18937_11636# ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1125 a_17695_15279# a_17507_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1126 a_8386_11247# net9 a_8217_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X1127 VGND a_12127_7093# uio_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1128 a_7929_7663# ts.o_res\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1129 a_11435_8864# _089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1131 a_8287_5487# a_7663_5493# a_8179_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1132 VGND a_7067_13812# _032_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1133 ts.ts_core.dac_vout_ana_ net14 a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1134 a_10229_9839# _066_ a_10147_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1135 a_8386_11247# net8 a_8300_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1136 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1137 a_1276_11293# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1138 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1139 VPWR clknet_2_2__leaf_clk a_855_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1140 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1141 VGND net69 a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1142 VPWR a_14287_4943# a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1144 VGND a_15483_1135# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1145 a_5922_8207# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1146 a_18293_4020# ui_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1147 VPWR a_16043_8359# a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
R14 uio_out[0] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1148 a_11812_5193# a_12547_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1149 a_7067_13812# _207_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1150 VPWR a_4135_11445# net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1151 a_10335_3029# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1152 a_8500_1929# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1153 a_3981_8449# a_3763_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1154 VGND a_11127_15797# a_11061_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1155 VGND _123_ a_11435_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X1156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1157 a_4349_17429# a_4131_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1158 VGND a_2111_11231# ts.ts_ctrl.temp_ctr\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1159 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1160 a_5043_13322# _210_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1161 a_12149_9295# ts.ts_ctrl.temp_ctr\[9\] a_11711_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1162 VPWR _143_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1163 a_16315_2223# a_16127_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1164 a_17599_6031# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
X1165 ts.ts_core.dac_vout_ana_ net14 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1166 a_6277_1455# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1167 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_17783_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1168 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1169 a_10154_5853# ts.ts_ctrl.temp_ctr\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1171 a_1633_7119# a_1589_7361# a_1467_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1173 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1174 VPWR a_11803_2767# a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1175 _114_ _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1176 ts.ts_core.dac_vout_ana_ net14 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1177 uio_out[5] a_14584_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X1178 a_11045_1367# a_11141_1109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1179 a_13560_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1180 _126_ a_10147_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1181 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9227_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1182 a_14475_5205# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1183 a_17143_7381# a_16955_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1184 _109_ a_11339_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X1185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1186 VPWR ts.ts_ctrl.state\[1\] _063_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1187 a_7719_17833# a_7203_17461# a_7624_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1188 VPWR a_7293_13077# a_7183_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1189 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1190 a_14384_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1191 a_16109_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1192 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1193 a_10980_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1194 ts.ts_core.dac_vout_ana_ net15 a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X1195 ts.ts_core.dac_vout_ana_ net14 a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1196 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1197 ts.ts_core.dac_vout_ana_ net72 a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1199 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1200 VPWR a_7313_4917# a_7343_5270# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1201 a_14852_8751# _108_ a_14584_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1202 a_16661_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X1203 a_7624_17821# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1205 a_6240_12711# ts.o_res\[8\] a_6382_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1206 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1207 VGND a_8399_18543# net8 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1208 a_17051_3029# a_16863_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1209 a_8657_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1210 a_6658_11293# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1211 a_16109_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1212 a_14015_10357# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X1213 a_13556_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1214 VGND net69 a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1215 a_4135_11231# a_3960_11305# a_4314_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1216 VGND net69 a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1217 a_13453_12381# _067_ a_13365_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1218 a_11969_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1219 VPWR a_15951_2919# a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1220 a_13046_4399# a_11969_4405# a_12884_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1221 a_2787_10205# ts.ts_ctrl.temp_ctr\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1223 VPWR a_15399_12711# a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1224 a_11991_1941# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1225 a_1761_3855# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1226 ts.ts_ctrl.temp_ctr\[16\] a_4503_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1227 a_1276_7119# _009_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1228 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.capload\[0\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1230 ts.ts_ctrl.temp_ctr\[1\] a_11035_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1231 a_1479_12925# a_855_12559# a_1371_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1232 a_3478_5487# a_2401_5493# a_3316_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1233 _055_ a_8235_8790# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1234 a_7105_1455# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1235 a_12591_6895# _062_ _114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1237 net15 a_11975_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1238 uo_out[7] a_9112_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1239 a_12792_15657# a_11877_15285# a_12445_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1240 ts.ts_core.dac_vout_ana_ net14 a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1241 VPWR a_7364_3855# a_7539_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1242 a_10378_15101# a_9301_14735# a_10216_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1243 a_8851_3285# a_8695_3553# a_8996_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X1244 a_11056_5193# _156_ a_10883_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1245 VPWR a_16403_10383# a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1246 a_6883_14887# ts.ts_ctrl.state\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1247 ts.ts_ctrl.temp_ctr\[13\] a_8459_17759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X1248 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _065_ a_16170_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R15 net32 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1249 a_5381_11225# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1250 a_4328_8207# a_3413_8207# a_3981_8449# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1251 ts.ts_core.dac_vout_ana_ net14 a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1252 _052_ a_9063_8534# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X1253 a_16569_10383# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1255 VPWR a_16043_7271# a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1256 a_8448_4007# ts.ts_ctrl.temp_ctr\[19\] a_8590_4182# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1257 a_9415_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 a_14664_12809# a_15399_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X1259 VGND net20 a_7337_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1260 VGND net69 a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1261 a_3576_12381# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1262 a_16569_1455# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1263 a_14296_4399# a_15031_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1264 a_12792_15657# a_11711_15285# a_12445_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1265 a_9267_18582# a_9085_18582# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1266 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1267 _039_ a_9871_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1268 VGND net68 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1269 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1270 a_5511_14735# a_5161_14735# a_5416_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1271 VPWR a_14663_5461# a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X1272 a_9500_12015# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1273 VPWR a_9112_11989# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1274 _066_ net10 a_16143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1275 _193_ ts.ts_ctrl.temp_ctr\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1276 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1277 VPWR _154_ a_9093_4438# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
R16 VGND net28 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1278 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1279 a_14545_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1280 VGND a_1459_14423# _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1281 a_9393_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1282 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1283 a_17673_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1284 VPWR _172_ a_4259_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1285 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1286 _159_ a_10294_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1287 a_10686_10383# ts.o_res\[0\] a_10605_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X1288 a_3825_15645# _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1289 a_12047_6835# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1290 VPWR a_6557_7637# a_6447_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1291 a_11159_6575# ts.ts_ctrl.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1292 a_9500_12015# ts.o_res\[15\] a_9112_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1293 a_15649_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1294 ts.ts_core.dac_vout_ana_ net71 a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1295 ts.ts_ctrl.temp_ctr\[6\] a_4411_12319# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1296 a_6741_4373# a_6523_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1297 a_6780_16911# _114_ a_6690_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X1298 a_3300_11293# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1299 VGND a_8877_15797# a_8811_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1300 ts.o_res\[14\] a_11127_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1301 a_3329_14985# ts.ts_ctrl.temp_ctr\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1302 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_16127_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1303 VPWR ts.o_res\[11\] a_10055_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X1304 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1305 VGND a_15465_3311# a_15571_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X1306 a_13731_8751# a_13551_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1307 VPWR a_8459_17759# ts.ts_ctrl.temp_ctr\[13\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1308 a_15465_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1309 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1310 VGND net68 a_16863_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1311 VPWR a_16495_10927# a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1312 a_10068_13423# _057_ a_9800_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1313 a_6704_3855# _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1314 a_17581_10159# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X1315 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1316 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1317 a_5043_13322# _210_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1318 VGND a_4871_17759# ts.ts_ctrl.temp_ctr\[11\] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1319 a_12993_4777# a_11803_4405# a_12884_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1320 VPWR a_10023_4917# a_10010_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1321 VGND net17 a_10557_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1322 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1323 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1324 a_3517_14569# a_2327_14197# a_3408_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1325 VGND net69 a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1326 a_8590_4182# _153_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1327 a_9414_3311# a_8656_3427# a_8851_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X1328 a_12218_3311# a_11141_3317# a_12056_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 a_17695_4399# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1330 VGND a_17783_5487# net14 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1331 a_14567_6575# a_14379_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1332 a_13859_13423# net12 a_13755_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X1333 ts.ts_core.dac_vout_ana_ net14 a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1334 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1335 a_14660_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1336 ts.o_res\[8\] a_5607_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1337 a_12243_15101# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1338 VPWR _143_ a_18969_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1339 a_9093_4438# ts.ts_ctrl.temp_ctr\[0\] a_8879_4438# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X1340 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1341 VGND a_5423_4917# net16 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1342 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1343 VGND a_10961_13799# _057_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1344 VPWR a_13919_3855# a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1345 a_1589_12801# a_1371_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1346 uo_out[4] a_9340_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1347 a_9256_11471# ts.o_res\[4\] a_9340_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1348 a_8761_12559# ts.ts_ctrl.temp_ctr\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1349 VGND _083_ a_8193_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1350 _019_ _183_ a_6185_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1351 a_9702_18365# a_9576_18267# a_9298_18251# VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1352 a_5455_6031# ts.ts_ctrl.temp_ctr\[18\] a_5361_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1353 _108_ a_12449_9301# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1354 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X1355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1356 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1357 a_8105_15285# a_7939_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1358 a_14567_6575# a_14379_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1359 a_16661_11247# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1360 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1362 VPWR _070_ a_11573_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1363 VGND net69 a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1364 a_12819_2223# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1365 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1366 a_15591_5487# ts.ts_ctrl.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1367 a_11285_10927# _052_ a_11456_11247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1368 uo_out[0] a_8836_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1369 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1370 _147_ a_11467_5825# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1371 a_16499_12821# a_16311_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1372 a_13556_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X1373 VPWR net67 a_16403_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1374 VPWR a_9195_15583# a_9182_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1375 VPWR a_12537_4373# a_12427_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
R17 VGND uio_out[1] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1376 net54 clknet_2_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1377 a_9629_13103# net8 a_9800_13423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1378 VPWR _114_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1379 VGND net5 a_17599_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1380 VGND net70 a_16955_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1381 a_12353_14977# a_12135_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1382 VPWR a_2969_5461# a_2859_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1383 a_17121_4943# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1384 VGND a_11272_11471# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1385 VPWR a_3583_14495# ts.ts_ctrl.temp_ctr\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1386 _176_ a_4259_14557# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1387 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13463_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X1388 VGND a_2375_12247# _167_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1389 a_7838_14191# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1390 a_12967_15583# a_12792_15657# a_13146_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1391 a_8933_4943# a_8767_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1392 VPWR a_12445_15253# a_12335_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1393 VPWR net68 a_17507_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1394 ts.ts_core.dac_vout_ana_ net71 a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1395 a_1371_9129# a_1021_8757# a_1276_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1396 a_16477_12559# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1397 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X1398 VPWR _074_ _094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X1399 VPWR clknet_2_3__leaf_clk a_9871_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1400 VPWR a_17507_15279# a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1401 VPWR a_9800_13423# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1402 ts.o_res\[11\] a_10299_16885# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1403 VGND clknet_2_2__leaf_clk a_855_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1404 a_10980_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1405 a_9669_9545# ts.ts_ctrl.temp_ctr\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1406 a_9209_16911# a_9043_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1407 a_16569_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1408 a_15212_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1410 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1411 VPWR _068_ a_14177_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X1412 VPWR clknet_0_clk a_4513_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1413 a_6699_12886# ts.o_res\[8\] a_6240_12711# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1414 a_3670_5853# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1415 VPWR a_5607_12533# a_5594_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1416 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1417 VPWR _062_ a_12357_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1418 a_15671_11733# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1419 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1420 a_11141_3317# a_10975_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1421 a_7026_4943# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1422 VPWR a_6076_14735# a_6251_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1423 VGND a_7365_15975# net66 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1424 a_2111_12533# a_1936_12559# a_2290_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1425 VPWR a_2397_15511# net64 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1426 a_5232_6005# _137_ a_5361_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1427 a_4515_4399# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1428 a_14475_6293# a_14287_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1429 a_11785_14735# a_11619_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1430 VGND a_6669_12533# a_6603_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1431 a_18763_8359# _139_ a_18937_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1432 VGND clknet_2_0__leaf_clk net53 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1433 VGND a_11207_7637# uio_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1434 VPWR net63 a_4798_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1435 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1436 VPWR a_16687_9447# a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1437 a_6879_11293# ts.ts_ctrl.temp_ctr\[7\] a_6516_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1438 a_15465_3311# a_15229_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X1439 a_11812_841# a_12547_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1440 a_15948_9295# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1441 VGND net68 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1442 VPWR a_3431_9839# _172_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1443 VPWR net69 a_17415_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1445 a_14545_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1446 VPWR a_16127_591# a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1447 ts.ts_core.dac_vout_ana_ net72 a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1448 VPWR a_12231_3615# ts.ts_ctrl.state\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1449 VPWR net67 a_11803_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1450 a_6523_9295# a_6173_9295# a_6428_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1451 VPWR a_11803_1679# a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1452 a_7737_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1454 a_11902_14557# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1455 VPWR a_7079_11445# a_7066_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1456 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1457 VGND clk a_7286_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1458 VGND ts.ts_core.dcdel_capnode_ana_ a_11057_591# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1459 VPWR net67 a_8491_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1460 a_12267_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1461 a_15308_7369# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1462 VPWR a_9227_1135# a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1464 a_10335_4117# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1465 VPWR a_9971_743# a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1466 a_2751_15253# ts.ts_ctrl.temp_ctr\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1467 VPWR a_14526_14165# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.135 ps=1.27 w=1 l=0.15
X1468 VPWR _093_ a_12181_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1469 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1470 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1471 ts.ts_ctrl.state\[1\] a_13059_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1472 a_1371_7119# a_855_7119# a_1276_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1473 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1474 VPWR a_14347_3615# ts.ts_ctrl.state\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1475 a_16661_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1476 a_5147_4703# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1477 a_1671_11471# ts.ts_ctrl.temp_ctr\[4\] _165_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1478 VGND a_18753_10548# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1479 a_7013_9129# a_5823_8757# a_6904_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1480 a_16591_1135# a_16403_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1481 VPWR a_4219_5461# _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X1482 ts.ts_core.dac_vout_ana_ net15 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1483 a_7364_3855# a_6283_3855# a_7017_4097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1484 _008_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1485 a_5989_11471# a_5823_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1486 a_11359_12015# net9 _051_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1487 a_13231_12247# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.141 ps=1.33 w=0.42 l=0.15
X1488 a_4259_14557# ts.ts_ctrl.temp_ctr\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1489 VPWR a_12547_4007# a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1490 a_10294_7093# ts.ts_ctrl.temp_ctr\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1491 a_8811_9295# ts.ts_ctrl.temp_ctr\[16\] a_8448_9447# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1492 a_14295_2919# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1493 _111_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1494 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X1495 a_14935_1941# a_14747_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1496 a_17051_1941# a_16863_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1497 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1498 a_14475_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1499 a_16591_10645# a_16403_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1500 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1501 VGND clknet_2_1__leaf_clk a_7663_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1502 a_14388_2223# a_15123_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1503 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1504 VPWR a_17507_15279# a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1505 a_17695_6575# a_17507_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1506 a_11767_17833# a_11417_17461# a_11672_17821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1507 a_12007_16150# ts.ts_ctrl.temp_ctr\[10\] a_12007_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1508 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1509 a_16209_9839# _099_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X1510 ts.ts_ctrl.state\[0\] a_12231_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1511 ts.ts_ctrl.state\[2\] a_14347_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1513 a_10202_4943# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1514 a_15741_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1515 a_15649_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1516 a_12952_13423# _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X1517 a_9232_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1518 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1519 a_10405_9545# ts.o_res\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1520 a_11812_4105# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1521 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1522 VPWR _140_ a_17877_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.117 ps=1.24 w=1 l=0.15
X1523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1524 a_12449_9301# _105_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1525 a_8877_15797# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1526 a_12997_6031# net5 a_12777_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X1527 ts.ts_ctrl.temp_ctr\[4\] a_2111_11231# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X1528 a_16499_12821# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1529 a_17121_4943# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1530 VPWR _069_ a_10975_8864# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1531 VPWR _067_ _094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1532 VGND _096_ a_11931_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1533 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1534 a_11785_14735# a_11619_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1535 ts.ts_core.capload\[13\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1536 a_17695_15279# a_17507_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1537 a_9339_18582# ts.o_res\[12\] a_9267_18582# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1538 a_7759_1135# a_7571_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1539 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1540 a_9301_14735# a_9135_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1541 VGND clknet_0_clk a_4986_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1542 a_6839_853# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1543 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1544 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1545 a_6631_9661# a_6007_9295# a_6523_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1546 a_8619_2223# a_7921_2229# a_8362_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
R18 VGND net25 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1547 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1549 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1550 VPWR a_12631_2223# a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1551 a_15741_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1552 a_18691_7663# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1553 VGND a_12777_6005# _144_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1554 a_6557_8725# a_6339_9129# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1555 a_3897_15645# _178_ a_3825_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1556 a_12007_15823# a_11753_16150# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1557 VPWR a_3613_10901# a_3503_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1558 a_15763_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1559 a_14461_11293# _073_ a_14355_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X1560 a_17603_9839# a_17415_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1561 a_3408_14569# a_2493_14197# a_3061_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1562 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1563 a_11808_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1564 a_4687_4917# a_4512_4943# a_4866_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1565 _128_ a_10975_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.26 ps=1.45 w=0.65 l=0.15
X1566 VGND a_8816_6183# _203_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1567 a_8816_6183# ts.ts_ctrl.temp_ctr\[1\] a_8958_6358# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1568 a_14063_10901# _074_ a_14461_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1569 VPWR a_12313_12234# net21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1570 ts.ts_ctrl.temp_ctr\[10\] a_4503_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1571 VGND net67 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1572 VPWR a_10294_7093# _159_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.135 ps=1.27 w=1 l=0.15
X1573 a_12489_15645# a_12445_15253# a_12323_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1574 VGND a_12047_6835# _061_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1575 VGND net69 a_16495_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1576 a_13183_7983# _113_ a_13601_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1577 a_17029_14735# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1579 VPWR a_18243_1135# net71 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1580 a_7013_8041# a_5823_7669# a_6904_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1581 a_7250_6575# a_6173_6581# a_7088_6953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1582 a_18836_12711# net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1583 a_12547_743# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1585 a_17581_10159# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1586 a_17143_7381# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1587 _156_ ts.ts_ctrl.state\[0\] a_9957_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1588 VGND net16 a_4669_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1589 uo_out[0] a_8836_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1590 a_15948_9295# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1591 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1592 a_4625_4373# a_4407_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1593 a_7263_4703# a_7088_4777# a_7442_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1594 a_9298_18251# a_9615_18141# a_9573_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1595 a_10321_9545# _106_ a_10239_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1596 VPWR ts.o_res\[9\] a_11285_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1597 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1598 uo_out[5] a_9524_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X1599 a_9440_12559# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1600 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_16311_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1601 VGND a_13546_10535# _090_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X1602 VPWR ts.ts_ctrl.temp_ctr\[8\] a_5271_13216# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1603 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1604 a_1936_11305# a_1021_10933# a_1589_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1605 a_13928_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1606 a_16591_10645# a_16403_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1607 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1608 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1609 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1610 VGND _159_ a_1855_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1611 a_12332_17833# a_11251_17461# a_11985_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1612 a_15212_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1613 a_14471_8207# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R19 VGND net30 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1614 VPWR ts.ts_ctrl.state\[2\] a_4075_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1615 VGND net69 a_15483_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1616 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1617 VPWR a_9227_1135# a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1618 a_11793_9545# _087_ a_11877_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1619 a_17143_8469# a_16955_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1620 a_8619_2223# a_7755_2229# a_8362_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1621 a_8907_16150# ts.o_res\[15\] a_8448_15975# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1622 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1623 a_6059_6005# _136_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X1624 a_13603_12533# net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X1625 a_8583_12559# _082_ a_8761_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1626 VGND _137_ a_5179_16367# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1627 ts.ts_core.dac_vout_ana_ net15 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1628 a_11902_14230# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1629 a_12085_12381# _072_ a_12013_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1630 VGND a_9524_12559# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1631 VGND _047_ a_9440_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X1632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1633 a_7183_13103# a_6559_13109# a_7075_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1634 VGND net16 a_7061_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1635 a_3933_12381# a_3889_11989# a_3767_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1636 net71 a_18243_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1637 VGND _075_ a_8745_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1638 a_9301_14735# a_9135_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1639 VPWR a_16403_10383# a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1641 a_5353_13469# ts.ts_ctrl.temp_ctr\[8\] a_5271_13216# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1642 ts.ts_core.dac_vout_ana_ net15 a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 VGND _182_ _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1644 _105_ a_11711_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1645 a_11969_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1646 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1647 a_12165_3689# a_10975_3317# a_12056_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1648 a_14281_3689# a_13091_3317# a_14172_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1649 VPWR _069_ _097_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1650 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1653 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1654 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1655 a_7026_6358# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1656 a_17695_15279# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1657 _059_ net11 a_14471_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1659 a_14901_13423# net12 a_15259_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VGND a_17332_3829# net67 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1661 a_13901_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1662 VPWR clknet_0_clk a_8022_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1663 ts.ts_core.capload\[12\].cap.Y net25 a_6185_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1664 a_9236_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1665 ts.ts_core.dac_vout_ana_ net47 a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1666 VPWR a_6629_15975# net58 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1667 ts.ts_core.dac_vout_ana_ net72 a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1668 a_7017_4097# a_6799_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1669 VPWR a_18763_9447# _152_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1670 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1671 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_18243_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1672 a_12797_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1673 a_14384_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1674 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 a_1769_7663# _138_ _160_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1676 a_8679_3029# a_8491_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1677 ts.ts_core.dac_vout_ana_ net72 a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1678 a_12135_14735# a_11785_14735# a_12040_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1679 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1680 ts.ts_ctrl.temp_ctr\[7\] a_4135_11231# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1681 a_7313_6005# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1682 a_4237_3855# a_3247_3855# a_4111_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1683 a_16609_6575# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1684 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1685 VGND net68 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1686 a_18937_11636# ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1687 a_8235_9117# a_7981_8790# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1688 VGND net69 a_17415_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1689 VGND net18 a_3657_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1690 a_9298_18251# a_9576_18267# a_9532_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1691 VGND _145_ a_15483_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1692 VGND net21 a_11597_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1693 a_6523_4777# a_6007_4405# a_6428_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1694 a_4407_4777# a_3891_4405# a_4312_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1695 VPWR a_16043_8359# a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X1696 VPWR _064_ a_14500_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1697 VGND a_3431_9839# _172_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1698 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1699 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16955_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1701 VPWR a_9615_18141# a_9576_18267# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1702 a_14471_13423# net11 _059_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1703 a_13560_841# a_14295_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1704 ts.ts_ctrl.temp_ctr\[11\] a_4871_17759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1705 a_3668_15823# _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1706 VGND a_6427_13621# _187_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1707 a_5607_14735# a_5161_14735# a_5511_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1708 a_16407_9839# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _100_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
X1709 a_3299_12533# _114_ a_3730_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X1710 VPWR a_5147_4703# a_5134_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1711 a_8836_10901# _048_ a_9224_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1712 a_15259_13423# net12 a_14901_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1713 _143_ _122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1714 a_12321_12705# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1715 _047_ net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1716 a_15321_7663# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X1717 a_16499_12821# a_16311_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1718 VGND net70 a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1719 a_14907_9545# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1720 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1722 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1723 a_13959_10429# a_13905_10535# a_13859_10429# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1724 VGND _067_ a_13445_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X1725 a_11587_3689# a_11141_3317# a_11491_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1726 a_13703_3689# a_13257_3317# a_13607_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1727 a_11760_14423# ts.ts_ctrl.temp_ctr\[9\] a_11902_14230# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1728 VPWR a_17783_5487# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1729 a_6858_16687# _188_ a_6563_16687# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X1730 VPWR a_11803_2767# a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1732 _114_ _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1733 ts.ts_core.dac_vout_ana_ net14 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1734 VGND a_18763_8359# _151_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1735 VPWR _177_ _178_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1736 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1737 VGND clknet_2_1__leaf_clk net55 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1738 a_11719_2197# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1740 a_13560_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1741 a_16315_853# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1742 VGND ts.ts_core.dac.vdac_single.en_pupd a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1743 VGND net69 a_16311_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1744 VGND net18 a_4025_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1745 a_17143_7381# a_16955_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1746 ts.ts_core.dac_vout_ana_ net14 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1747 VPWR a_18234_10927# net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1748 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1749 a_4535_14557# ts.ts_ctrl.temp_ctr\[10\] a_4429_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1750 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1751 VGND a_2014_3967# a_1972_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1752 a_7847_7663# _090_ a_7929_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1753 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1754 a_7286_9839# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1755 a_4131_17833# a_3781_17461# a_4036_17821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1756 a_5085_5487# net59 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1757 a_9340_11471# _051_ a_9608_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1758 a_16960_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1759 VPWR a_12789_13077# _101_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X1760 VGND net20 a_8399_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1761 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1762 a_14445_9545# _135_ a_14717_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1763 VPWR _059_ a_16187_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1764 VGND ts.ts_core.dac.vdac_single.en_pupd a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1765 VPWR a_16311_12559# a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1766 VGND _177_ a_4713_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X1767 a_11272_11471# ts.o_res\[10\] a_11188_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1768 a_8287_5487# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1769 VPWR a_6741_6549# a_6631_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1770 VPWR clknet_2_1__leaf_clk a_9779_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1771 ts.ts_core.dac_vout_ana_ net72 a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1772 a_17143_8469# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1773 a_17695_8751# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 VGND a_5179_16367# _138_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1776 a_14660_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1777 VGND _211_ a_12228_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X1778 a_12127_7093# a_12493_7369# a_12851_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1779 ts.ts_core.capload\[0\].cap.Y net22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1780 VPWR net12 a_15451_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1781 a_13923_1135# a_13735_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1783 a_12752_12809# _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1784 VPWR a_10513_6273# a_10403_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1785 a_17051_3029# a_16863_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1786 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1787 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1788 VPWR a_6884_5095# _221_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1789 uo_out[2] a_11272_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1791 a_7026_5270# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1792 a_3960_11305# a_3045_10933# a_3613_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1793 a_11969_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1794 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1795 a_1846_4221# a_1573_3855# a_1761_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1796 _099_ _065_ a_14189_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1797 a_17695_8751# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1798 ts.ts_core.dac_vout_ana_ net14 a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X1799 VPWR a_8399_18543# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1800 a_11808_3855# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1801 a_4036_17821# _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1802 a_17695_15279# a_17507_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1803 a_17143_8469# a_16955_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1804 uo_out[6] a_9800_13423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1805 VPWR ts.o_res\[6\] a_9629_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1806 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1807 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1808 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1809 a_2045_12559# a_855_12559# a_1936_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1810 VPWR a_16587_7663# a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1812 VPWR _138_ a_3413_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1813 VGND _073_ a_15159_11248# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1815 a_7929_7983# ts.ts_ctrl.temp_ctr\[19\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1816 ts.ts_core.dac_vout_ana_ net14 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1817 a_9865_7369# _158_ a_9781_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1818 a_17121_7119# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1819 a_14259_11293# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X1820 a_3762_14557# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1821 a_14567_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1822 VPWR a_16043_7271# a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X1823 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1824 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1826 net69 a_18234_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1827 a_13042_13423# _072_ a_12952_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1828 a_7013_11471# a_5823_11471# a_6904_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1829 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1830 a_12591_11159# ts.ts_core.o_tempdelay VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X1831 a_9297_13423# ts.o_res\[12\] a_8859_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1832 a_11977_13423# ts.ts_ctrl.temp_ctr\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1833 VPWR a_8787_2197# a_8703_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1834 a_16170_6895# _065_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1835 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1836 a_14545_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1838 a_13556_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1839 a_8807_4438# a_8625_4438# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1840 _102_ a_11895_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1841 VPWR a_3944_14709# _179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1842 a_9393_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1843 VPWR a_18847_14709# net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1845 a_11991_1941# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1846 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1847 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10147_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1848 a_10975_9295# _126_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X1849 VGND _061_ a_13992_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.0662 ps=0.735 w=0.42 l=0.15
X1850 a_7285_12015# ts.ts_ctrl.temp_ctr\[11\] a_7203_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1851 a_2843_14569# a_2493_14197# a_2748_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1852 a_11808_3855# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1853 a_9960_9071# ts.ts_ctrl.state\[0\] a_9770_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X1854 ts.ts_core.dac_vout_ana_ net71 a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1855 VGND _144_ a_8241_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1856 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1857 a_12335_15279# a_11711_15285# a_12227_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1858 VPWR a_2271_4221# a_2439_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1859 VGND net18 a_5037_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1860 a_7066_11837# a_5989_11471# a_6904_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1862 a_6173_9295# a_6007_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1863 a_17699_13799# net69 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1864 a_18937_2932# ui_in[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1866 a_3663_15511# _114_ a_3897_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1868 a_10335_3029# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1869 a_8500_1929# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1870 a_9681_9295# ts.o_res\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1872 VPWR a_12700_14735# a_12875_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1873 a_2787_10205# _162_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1874 _083_ a_14526_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X1875 a_2537_9323# _159_ a_2451_9323# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1876 a_16315_2223# a_16127_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1877 VGND ts.ts_ctrl.state\[1\] a_12596_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1878 a_8877_15797# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1879 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1880 VGND a_11045_1367# net57 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1881 VPWR _187_ _188_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1882 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1883 VGND a_6792_7271# _204_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1884 a_11812_5193# a_12547_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X1885 ts.ts_core.capload\[2\].cap.Y net30 a_5909_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1886 VGND net68 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X1887 a_6541_17999# a_6375_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1888 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R20 ts.ts_core.capload\[13\].cap_26.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1889 a_10299_16885# a_10124_16911# a_10478_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1890 a_16589_5193# net6 a_16465_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.235 ps=1.47 w=1 l=0.15
X1891 a_17143_7381# a_16955_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X1892 a_13832_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1893 VPWR _215_ a_9871_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1895 VPWR _081_ a_8749_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1896 a_14024_8207# _065_ a_13834_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1897 VPWR a_16403_10383# a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1898 VPWR _143_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1899 a_2873_12335# _168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1900 VGND a_17783_5487# net14 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1901 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1902 a_1633_11293# a_1589_10901# a_1467_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1903 a_6725_13109# a_6559_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1904 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1905 a_14384_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1906 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1907 a_17029_2767# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1908 VPWR a_13919_3855# a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X1909 VGND a_2659_10357# a_2401_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X1910 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1911 ts.ts_core.dac_vout_ana_ net72 a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1912 a_6785_9295# a_6741_9537# a_6619_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1913 a_12007_16150# ts.o_res\[10\] a_11935_16150# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1914 VGND net67 a_6651_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1915 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1916 a_8856_10383# ts.o_res\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1917 VPWR _195_ a_3479_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1918 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1919 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1920 a_17051_3029# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1921 VGND net17 a_8441_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1922 a_16170_6895# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1923 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1924 _132_ a_8583_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X1925 VPWR _172_ a_4126_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X1926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1927 a_11969_4405# a_11803_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1928 a_8919_5791# a_8744_5865# a_9098_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1929 a_2290_9117# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1930 VPWR a_4696_17833# a_4871_17759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1931 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1932 VPWR a_11207_7637# uio_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1933 VGND _083_ a_7549_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1934 a_14384_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1935 VPWR a_8877_15797# a_8907_16150# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1936 a_10441_5785# ts.ts_ctrl.temp_ctr\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1937 a_16109_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1938 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1939 _094_ _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X1940 VGND net18 a_1633_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1941 _145_ a_8155_4737# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1942 VGND a_10018_4373# a_9976_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1943 _065_ _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1944 a_11851_12247# ts.o_res\[10\] a_12085_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1945 net15 a_11975_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1946 VGND clknet_2_3__leaf_clk a_9135_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1947 a_6557_8725# a_6339_9129# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1948 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1949 VPWR net6 a_15321_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1951 ts.o_res\[3\] a_7079_9055# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1952 a_17029_14735# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1953 _170_ ts.ts_ctrl.temp_ctr\[7\] a_2695_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1954 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
R21 VPWR ts.ts_core.capload\[8\].cap_36.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1956 a_16683_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1957 a_3408_14569# a_2327_14197# a_3061_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1958 VPWR a_6983_15797# a_6725_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X1959 a_6833_15253# a_6615_15657# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1960 a_7355_15583# a_7180_15657# a_7534_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1962 a_13611_4917# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1963 a_7815_17833# a_7369_17461# a_7719_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1964 VGND a_4279_4123# a_4237_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1965 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_17332_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1966 a_8447_6196# _203_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1968 _004_ a_11056_5193# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
X1969 VPWR ts.ts_ctrl.temp_ctr\[6\] a_2695_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1970 a_6428_9295# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1971 a_10387_15823# a_9871_15823# a_10292_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1972 a_10980_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1973 VPWR a_2111_12533# a_2098_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1974 a_5786_12559# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1975 VGND clknet_2_0__leaf_clk a_2235_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1976 VGND _134_ a_14195_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1977 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1978 a_10417_9295# ts.o_res\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1979 a_6516_11159# ts.o_res\[7\] a_6658_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1981 a_16109_6031# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1982 a_1858_12335# _164_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X1983 a_15763_4117# a_15575_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1984 a_9063_8534# ts.o_res\[17\] a_8991_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1985 a_13556_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1986 a_17673_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1987 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1988 VPWR a_12547_743# a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1989 VPWR a_16311_12559# a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1991 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1992 a_11285_10927# ts.o_res\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1993 a_7937_17429# a_7719_17833# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1994 uio_out[6] a_12127_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1995 VPWR a_14663_5461# a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X1996 a_14660_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1997 ts.ts_core.dac_vout_ana_ net15 a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1999 a_3321_12021# a_3155_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2000 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2001 a_14015_10357# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X2002 a_3601_3855# net56 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2005 a_17673_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2006 a_8193_12335# ts.ts_ctrl.temp_ctr\[4\] a_7847_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2007 a_7526_4221# a_6449_3855# a_7364_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2008 a_9063_8207# a_8809_8534# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X2009 a_12221_16150# ts.ts_ctrl.temp_ctr\[10\] a_12007_16150# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X2010 a_12700_14735# a_11785_14735# a_12353_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2011 net68 a_13611_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2012 a_9669_9545# ts.o_res\[4\] a_9585_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2013 a_9236_841# a_9971_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2014 VPWR a_3408_14569# a_3583_14495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2015 VGND a_5607_12533# a_5541_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2016 a_17143_5205# a_16955_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2017 VGND net69 a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2018 a_10313_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2019 a_7247_6031# ts.ts_ctrl.temp_ctr\[17\] a_6884_6183# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2020 VPWR a_16495_12015# a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X2021 a_9440_12559# ts.o_res\[5\] a_9524_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2022 a_7369_17461# a_7203_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2023 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X2024 a_16569_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2025 _107_ a_10239_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2026 a_6904_9129# a_5823_8757# a_6557_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2027 VGND clknet_2_3__leaf_clk a_9043_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2028 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2029 VPWR clknet_2_3__leaf_clk a_9135_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2030 a_12267_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2031 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref _146_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2032 a_2847_5865# a_2401_5493# a_2751_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2033 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2035 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2036 a_1941_4221# a_1407_3855# a_1846_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2037 a_9792_12559# _056_ a_9524_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2038 a_16043_8359# ts.ts_core.dac.vdac_single.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2039 VGND net67 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2040 a_11207_7637# _096_ a_12181_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2041 a_4345_12393# a_3155_12021# a_4236_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2042 VPWR a_6247_17429# a_5989_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X2043 a_12040_14735# _036_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2044 VPWR a_10952_15823# a_11127_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2045 VPWR a_10147_1679# a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2046 a_3889_11989# a_3671_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2048 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2049 a_9415_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2050 ts.ts_ctrl.temp_ctr\[2\] a_2111_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X2051 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2052 _074_ a_17191_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2053 a_6515_10058# _219_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2054 a_2777_12559# ts.ts_ctrl.temp_ctr\[4\] a_2695_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2055 a_16591_1135# a_16403_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2056 a_17673_6895# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2057 ts.ts_core.dac_vout_ana_ net14 a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X2058 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2059 VPWR a_12547_4007# a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X2060 VPWR a_13919_3855# a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2061 ts.ts_ctrl.temp_ctr\[18\] a_4687_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2062 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2063 _138_ a_5179_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
R22 VPWR ts.ts_core.capload\[9\].cap_37.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2064 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2065 a_16683_12015# a_16495_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2066 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2067 VGND a_14707_10901# _075_ VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=1 as=0.0991 ps=0.955 w=0.65 l=0.15
X2068 a_18937_2932# ui_in[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2069 a_17051_1941# a_16863_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2070 a_1854_6575# _159_ a_1551_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X2071 a_1589_14977# a_1371_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2072 a_14545_6895# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2073 a_6904_11471# a_5989_11471# a_6557_11713# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2074 VPWR a_15299_13647# a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2075 VPWR a_7631_17973# ts.ts_ctrl.temp_ctr\[12\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2076 a_9061_16665# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2077 a_4503_15797# a_4328_15823# a_4682_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2078 _154_ a_9287_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2079 VGND _139_ a_11553_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2080 a_2111_11231# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2081 _062_ ts.ts_ctrl.state\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2082 a_17695_6575# a_17507_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2083 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2084 a_11207_7637# a_11573_7663# a_11931_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2085 VPWR net69 a_16495_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2086 a_1936_9129# a_1021_8757# a_1589_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2087 a_17143_14191# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2088 a_13599_6807# a_13963_6896# a_13921_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2089 VPWR a_3061_14165# a_2951_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2090 VGND a_3491_5791# ts.ts_ctrl.temp_ctr\[17\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2091 a_5989_8757# a_5823_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2092 a_13967_12711# net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
R23 ts.ts_core.capload\[12\].cap_25.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2093 VPWR a_15943_6031# a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2094 VGND _157_ _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2095 a_16043_7271# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2097 _172_ a_3431_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2098 VPWR _113_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2099 ts.ts_core.dac_vout_ana_ net15 a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2100 a_6244_11471# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2101 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2102 a_7355_15583# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2103 a_14901_13423# net12 a_15259_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2104 VPWR _211_ a_12221_16150# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
R24 tt_um_hpretl_tt06_tempsens_44.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2106 a_16315_5487# a_16127_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2107 VPWR a_12275_6281# _113_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2108 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2109 a_15487_13909# a_15299_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2110 VPWR a_12631_2223# a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X2111 a_13705_6353# _059_ a_13633_6353# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0441 ps=0.63 w=0.42 l=0.15
X2112 a_12313_12234# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2113 ts.ts_core.dac_vout_ana_ net72 a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2114 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2115 a_7759_1135# a_7571_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2116 a_9224_10927# ts.o_res\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2117 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2118 a_8193_7983# ts.o_res\[19\] a_7847_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2119 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd _065_ a_17599_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2120 VPWR a_2397_6807# net61 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2121 a_14663_5461# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2122 VPWR a_18234_10927# net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2123 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2124 a_11808_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2125 VGND _194_ a_4229_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2126 a_14296_4399# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2127 a_14986_9849# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.169 ps=1.5 w=0.42 l=0.15
X2128 VPWR a_12189_14489# a_12219_14230# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2129 VPWR _178_ a_3663_15511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2130 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X2131 VPWR a_15159_11248# a_14707_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X2132 VPWR a_12631_2223# a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2133 a_14475_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2134 VGND _097_ a_14418_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2135 a_1371_11305# a_855_10933# a_1276_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2136 _118_ a_10239_13897# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2137 a_16293_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2138 a_2751_6549# ts.ts_ctrl.temp_ctr\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2139 a_8448_9447# ts.ts_ctrl.temp_ctr\[16\] a_8590_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
R25 VGND uio_oe[2] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2140 _058_ a_12596_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2142 VPWR a_4135_11231# a_4122_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2143 a_9608_11471# ts.o_res\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2144 VPWR _214_ a_8767_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2145 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2146 a_17603_9839# a_17415_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2148 a_11188_11471# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2149 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2151 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_13183_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2152 a_16127_10159# _094_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2153 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2154 VPWR clknet_2_2__leaf_clk a_3155_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2155 VGND ts.ts_core.dcdel_capnode_ana_ a_9033_591# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2156 VPWR a_17935_13363# net70 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2157 a_12493_7369# _110_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2158 a_13183_7983# _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2159 a_11540_11471# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2160 VPWR net72 a_18243_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2161 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2162 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2163 a_12157_9813# _066_ a_12403_10177# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2164 a_10441_15577# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2165 ts.ts_core.dac_vout_ana_ net72 a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2166 a_14567_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2167 VPWR a_8399_18543# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2168 VPWR a_9643_14410# _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2169 a_17121_4943# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2170 a_6817_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2171 VPWR _080_ a_11131_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2172 VPWR a_16955_14191# a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2173 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2174 a_8500_1929# a_9235_1831# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2175 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2176 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2177 a_11812_5193# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2178 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2179 VGND _083_ a_12241_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2180 a_5081_17161# _137_ _181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2181 net19 a_8399_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2182 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2183 _042_ a_8031_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2184 a_13928_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2185 a_12013_12381# _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2187 a_8612_3311# a_8175_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2188 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2190 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2191 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2192 ts.ts_core.capload\[12\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2193 a_11753_3677# a_11709_3285# a_11587_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2194 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2195 a_15212_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2196 VGND _050_ a_11540_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X2197 a_14928_11293# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.104 ps=1 w=0.42 l=0.15
X2198 a_13836_11721# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2199 a_16683_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2200 a_18691_7663# _094_ _096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2201 a_5515_10357# a_5340_10383# a_5694_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2202 a_7473_3855# a_6283_3855# a_7364_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2203 a_12267_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2204 _134_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2205 a_4411_12319# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2206 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2207 a_11793_9545# _104_ a_11711_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2208 VPWR a_6427_16341# _021_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2209 ts.ts_core.dac_vout_ana_ net72 a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2210 ts.ts_core.dac_vout_ana_ net15 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2211 a_4165_5185# a_3947_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2212 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2213 VGND a_8787_2197# a_8745_2601# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2214 _140_ a_13643_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2215 a_6435_9129# a_5989_8757# a_6339_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2216 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2217 VPWR a_8448_9447# _219_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2218 a_8590_9622# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2220 VPWR ts.ts_ctrl.temp_ctr\[9\] a_4073_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2221 VPWR a_16180_11989# _067_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2222 a_14935_1941# a_14747_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2223 a_17051_1941# a_16863_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2224 VPWR _094_ a_15749_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2225 a_8163_8790# a_7981_8790# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2226 net13 a_18847_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2227 VGND a_6945_11225# a_6879_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2228 VPWR a_2751_6549# a_2493_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X2229 a_4680_11445# res2_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2230 ts.ts_core.dac_vout_ana_ net15 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2231 _140_ _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2232 _213_ a_12007_16150# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X2233 VPWR _138_ a_14907_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2234 ts.ts_core.dac_vout_ana_ net71 a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2235 a_6523_9295# a_6007_9295# a_6428_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2236 VGND _192_ a_4799_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X2237 a_3889_11989# a_3671_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2238 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2239 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2240 net19 a_8399_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2241 a_13901_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2242 VPWR _065_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X2243 a_11396_3677# _004_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2244 a_13512_3677# _006_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2245 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2246 VPWR a_14295_743# a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2247 VGND _094_ a_18243_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
X2248 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2249 VGND net8 a_8532_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2250 VGND res2_n a_6559_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2251 VPWR a_17507_4399# a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2252 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2253 VPWR a_3413_3311# a_3519_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X2254 a_6629_15975# a_6725_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X2255 a_13257_3317# a_13091_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2256 a_6895_3855# a_6449_3855# a_6799_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2257 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2258 VGND net68 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2259 a_16465_5193# net6 a_16311_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2260 VGND net9 a_7981_8790# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X2261 a_14584_8751# _097_ a_14500_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2262 _020_ a_6690_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2263 VPWR a_12884_4777# a_13059_4703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2264 VGND clknet_2_3__leaf_clk a_6375_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2265 VPWR ts.ts_ctrl.temp_ctr\[2\] a_1769_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X2266 a_1589_8725# a_1371_9129# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2267 a_4025_15823# a_3981_16065# a_3859_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2268 VPWR a_16863_14735# a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2269 _143_ _059_ a_13601_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2270 ts.ts_ctrl.temp_ctr\[3\] a_2111_9055# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2271 ts.ts_core.dac_vout_ana_ net14 a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X2272 _036_ a_11343_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2273 a_10275_4399# a_9411_4405# a_10018_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2274 VPWR net4 a_16609_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2275 VGND a_4871_17759# a_4805_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2276 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2277 VGND a_8468_10357# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2278 VPWR a_15399_12711# a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2279 VPWR a_14571_11623# a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X2280 VGND ts.ts_ctrl.state\[1\] a_13821_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2281 a_7197_6953# a_6007_6581# a_7088_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2282 VGND clknet_0_clk a_4986_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2283 VPWR a_6240_12711# _210_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2285 _106_ a_8491_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2286 ts.ts_ctrl.temp_ctr\[14\] a_7355_15583# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2287 a_4314_11293# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2288 net72 a_18335_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2289 a_16315_853# a_16127_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2290 a_1551_6807# _160_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X2291 a_12257_8457# _121_ a_12161_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2292 a_10686_10383# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X2293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2294 VGND _054_ a_8856_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2295 a_4236_12393# a_3321_12021# a_3889_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2296 a_4684_5487# _198_ a_4219_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X2297 a_6435_8041# a_5989_7669# a_6339_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2298 a_16683_12015# a_16495_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2299 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2300 a_6884_5095# ts.o_res\[18\] a_7026_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2301 a_14707_10901# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X2302 a_11057_591# net24 ts.ts_core.capload\[11\].cap.Y VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2303 _142_ a_18735_6059# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X2304 a_16569_10383# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2305 VGND a_8877_3829# a_8811_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2306 VPWR a_10147_2767# a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2307 VPWR _074_ a_12853_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X2308 a_8573_7663# ts.ts_ctrl.temp_ctr\[17\] a_8491_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2309 a_8500_1929# a_9235_1831# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X2310 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2311 a_17695_8751# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2312 a_4588_14709# _176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2313 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2314 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2315 VGND _061_ a_17599_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2316 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2317 a_4680_11445# res2_n VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2318 a_13923_1135# a_13735_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2319 a_5893_5719# a_5989_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X2320 VPWR clk a_7286_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2321 VPWR net11 a_16143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2322 a_17051_3029# a_16863_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2323 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2324 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2325 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2326 a_17029_14735# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2327 ts.ts_core.dac_vout_ana_ net14 a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2328 VGND clknet_0_clk a_4513_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2329 VGND a_4135_11231# a_4069_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2330 VGND _214_ a_8767_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2331 a_15487_13909# a_15299_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2332 a_2849_12559# ts.ts_ctrl.temp_ctr\[5\] a_2777_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
R26 ts.ts_core.capload\[6\].cap_34.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2333 a_12267_1135# a_12079_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2334 a_11812_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2335 ts.o_res\[7\] a_7079_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2336 VPWR a_13769_6296# a_13705_6353# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.0672 ps=0.74 w=0.42 l=0.15
X2337 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2338 a_6619_6953# a_6173_6581# a_6523_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2339 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_16863_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2340 _150_ a_17017_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.373 ps=1.75 w=1 l=0.15
X2341 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2342 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_13735_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2343 a_2098_12925# a_1021_12559# a_1936_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2344 a_14584_8751# _108_ a_14852_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2345 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2346 VPWR a_14295_2919# a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2347 a_14195_9545# _134_ a_14445_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2348 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2349 a_1936_9129# a_855_8757# a_1589_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2350 a_2355_4221# a_1573_3855# a_2271_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2352 a_16293_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2353 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2354 a_10229_9839# ts.o_res\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2355 VGND _027_ a_9414_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2356 VGND a_2755_8983# _162_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2357 VPWR a_18847_16341# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2358 a_1585_11721# _138_ _165_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2359 a_3730_12559# _169_ a_3435_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2360 a_9391_5309# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2361 a_1371_14735# a_1021_14735# a_1276_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2362 a_2397_6807# a_2493_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X2363 VGND a_9340_11471# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2364 a_9340_11471# ts.o_res\[4\] a_9256_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2365 _042_ a_8031_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2366 a_10471_5526# _112_ a_10012_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2367 a_2045_14191# _138_ _175_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2368 VGND a_16187_7895# _060_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2369 a_10321_13897# ts.ts_ctrl.temp_ctr\[14\] a_10239_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2370 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2371 VGND net69 a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2372 a_13859_10429# _067_ a_13755_10429# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X2373 a_6839_853# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2374 a_14545_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2375 a_4025_8207# a_3981_8449# a_3859_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2376 a_9559_16911# a_9043_16911# a_9464_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2377 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2378 VPWR a_10012_15511# _217_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2379 a_13546_13335# a_14015_13077# a_13959_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X2380 VPWR net17 a_8175_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2381 a_13079_6281# _140_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X2382 VGND net4 a_16170_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X2383 a_15649_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R27 VGND net35 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2384 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2385 VPWR a_6904_9129# a_7079_9055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2386 a_6723_15279# a_6099_15285# a_6615_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2387 VGND a_15483_1135# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2388 a_6601_8029# a_6557_7637# a_6435_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2389 VPWR ts.ts_ctrl.state\[2\] a_10975_8864# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2390 VGND _143_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2391 a_9245_6005# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2392 a_16293_13423# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2393 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2394 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2395 VPWR _059_ a_11437_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2396 VGND net69 a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2397 a_4437_15823# a_3247_15823# a_4328_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2398 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2399 a_6247_17429# ts.ts_ctrl.temp_ctr\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2400 VPWR a_2111_14709# ts.ts_ctrl.temp_ctr\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2401 a_8679_3029# a_8491_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2402 a_13836_11721# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2403 VPWR a_7719_15797# a_7461_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X2404 a_11285_10927# _050_ a_11456_11247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2405 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2406 a_9524_12559# _056_ a_9792_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2407 VPWR a_9227_2223# a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2408 a_11127_15797# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2409 a_16315_2223# a_16127_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2410 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2411 a_6515_5108# _221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2412 VGND net70 a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2413 ts.ts_core.dac_vout_ana_ net72 a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2415 ts.ts_core.dac_vout_ana_ net15 a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2416 a_16591_1135# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2417 a_7159_16599# ts.ts_ctrl.temp_ctr\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2418 a_2969_5461# a_2751_5865# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2419 a_12883_7983# _113_ a_12787_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.107 ps=0.98 w=0.65 l=0.15
X2420 a_18847_16341# uio_in[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2422 a_17673_9071# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2423 a_1677_14511# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2424 _007_ _157_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2425 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2426 a_10229_10159# _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2427 a_17051_3029# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2428 VGND net8 _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R28 VPWR tt_um_hpretl_tt06_tempsens_43.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2429 a_16315_13103# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2430 ts.ts_ctrl.temp_ctr\[12\] a_7631_17973# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X2431 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2432 _191_ a_5271_13216# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2433 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2434 a_14453_10205# ts.ts_core.i_precharge_n a_14353_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X2435 a_16477_12559# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2436 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2437 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2438 ts.ts_core.capload\[1\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2439 a_14384_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2440 a_6945_11225# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2441 a_6251_14709# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2442 a_6244_11471# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2443 _114_ _112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2444 VPWR a_10443_4373# a_10359_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2445 VGND ts.ts_core.dac.vdac_single.en_pupd a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2446 a_13146_15645# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2447 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2448 a_2045_9129# a_855_8757# a_1936_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2449 a_7718_3855# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2450 VPWR a_11119_4373# _005_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2451 VGND a_10012_5719# _157_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2452 ts.ts_core.dac_vout_ana_ net72 a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2453 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17599_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2454 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2455 a_15465_13647# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2456 a_17051_3029# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2457 a_5515_10357# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
R29 net36 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2458 a_7286_9839# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2459 a_13923_1135# a_13735_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2460 net56 a_3519_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2461 VGND _215_ a_9871_17455# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2462 a_9553_18582# ts.ts_ctrl.temp_ctr\[12\] a_9339_18582# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X2463 a_14901_13423# net10 a_14471_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X2464 VPWR a_17332_3829# net67 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2465 a_17051_3029# a_16863_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2467 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2468 a_6669_12533# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2469 _036_ a_11343_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2470 a_16109_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2471 VGND net69 a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2472 a_9161_3677# a_8782_3311# a_9089_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2474 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2475 VPWR a_18234_10927# net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2477 a_17143_8469# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2478 a_15671_11733# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2479 a_6244_9117# _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2480 VGND _061_ a_16170_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2481 VPWR _047_ a_9224_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X2482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2483 a_7759_1135# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2484 VPWR a_14287_4943# a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2485 a_12591_6895# _062_ _114_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2487 VPWR a_13599_6807# _115_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2489 a_8496_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2490 VPWR _066_ a_9687_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X2491 a_2951_14191# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2492 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2494 a_1479_7485# a_855_7119# a_1371_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2495 a_6669_12533# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2497 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2498 VGND _172_ a_4535_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2500 VPWR _172_ a_4713_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X2501 a_2290_12559# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2502 a_10335_4117# a_10147_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2503 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2504 a_14545_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2505 a_18787_12809# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.27 ps=2.54 w=1 l=0.15
X2506 a_3307_13799# _172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X2507 a_4798_17161# _177_ a_4495_16885# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X2508 VPWR _039_ a_10334_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2509 _051_ net9 a_11359_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2510 a_17603_9839# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2511 VGND net69 a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2512 a_10980_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2513 ts.ts_core.dac_vout_ana_ net47 a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2514 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16127_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X2515 a_4069_11305# a_2879_10933# a_3960_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2516 _010_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2517 a_1467_9129# a_1021_8757# a_1371_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2518 VGND ts.ts_core.dcdel_capnode_ana_ a_6181_591# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2519 a_4073_14985# _172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2520 VGND ts.ts_ctrl.state\[2\] _062_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2521 a_3316_5865# a_2235_5493# a_2969_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2522 a_8447_6196# _203_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2523 VGND _133_ a_14195_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2524 VPWR a_18937_2932# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2525 a_13560_841# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2526 a_17121_7119# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2527 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2528 VPWR a_13611_4917# net68 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2529 a_5449_10383# a_4259_10383# a_5340_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2530 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2531 a_5081_17161# _177_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2532 VPWR a_4503_15797# a_4490_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2533 a_14545_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2534 a_17143_14191# a_16955_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2535 a_11969_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2536 VPWR net67 a_16127_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2537 a_6247_5461# ts.ts_ctrl.temp_ctr\[18\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2538 VPWR a_1936_14735# a_2111_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2539 a_13556_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2540 a_9393_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2541 a_2656_5853# _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2542 a_17673_6895# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2543 VGND a_13603_12533# _068_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2544 VPWR a_4952_11159# _206_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2545 a_11359_12015# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2546 a_3686_4221# a_3413_3855# a_3601_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2547 VGND _159_ a_1769_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2548 ts.ts_core.dac_vout_ana_ net71 a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2549 VPWR _211_ a_9553_18582# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2550 VPWR a_16403_1135# a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2551 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2552 a_8657_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2553 a_4407_4777# a_4057_4405# a_4312_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2554 ts.ts_ctrl.temp_ctr\[8\] a_3583_14495# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X2555 VGND a_2111_12533# a_2045_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2556 a_11889_9295# ts.ts_ctrl.temp_ctr\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X2557 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2558 a_9393_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2559 VPWR net67 a_14379_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2560 a_11540_11471# _053_ a_11272_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2561 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2562 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2563 a_4883_10749# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2564 VPWR a_17507_15279# a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2565 a_11991_1941# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2566 VGND _058_ a_11053_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2567 a_14355_11293# _067_ a_14259_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X2568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2569 a_12507_17759# a_12332_17833# a_12686_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2570 a_9602_13974# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2571 VPWR a_11985_17429# a_11875_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2572 a_13556_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2573 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2574 a_17143_5205# a_16955_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2575 a_11808_4943# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2576 a_10313_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2577 a_17191_11445# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X2578 a_7549_12335# ts.ts_ctrl.temp_ctr\[7\] a_7203_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2579 ts.ts_core.dac_vout_ana_ net14 a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2580 a_4683_13077# ts.ts_ctrl.temp_ctr\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2581 VPWR a_18671_14451# net9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2582 a_4588_14709# _176_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2583 a_8906_5487# a_7829_5493# a_8744_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2584 VGND _081_ a_9297_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2585 ts.ts_ctrl.temp_ctr\[17\] a_3491_5791# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X2586 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2587 uio_out[4] a_11207_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2588 a_18937_8235# _150_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2589 a_16499_12821# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2590 a_14787_13693# a_14733_13799# a_14687_13693# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2591 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2592 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2593 a_15952_9545# a_16687_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2594 a_5729_14977# a_5511_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2595 a_17017_4399# _098_ a_16945_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X2596 VPWR a_11573_7663# a_11207_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2597 a_13086_11159# a_13555_10901# a_13499_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X2598 a_9602_13647# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X2599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2600 VPWR a_10147_1679# a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2601 _094_ _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=2.8 w=1 l=0.15
X2602 a_9415_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2603 VGND a_17783_5487# net14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2604 a_14545_6895# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2606 a_11343_12809# _118_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2607 a_5871_13335# _187_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2608 a_4687_4917# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2609 VGND net68 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2610 VPWR a_7571_1135# a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2611 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2612 VGND _183_ a_6880_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X2613 a_12700_14735# a_11619_14735# a_12353_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2614 VPWR a_13919_3855# a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2615 a_13086_11159# a_13445_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2616 VGND net67 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2617 net52 clknet_2_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2618 a_9651_14735# a_9301_14735# a_9556_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2619 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2620 a_7838_14191# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2621 VGND ts.ts_ctrl.state\[0\] a_11429_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2622 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2623 VPWR _128_ a_9751_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2624 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2625 a_4503_8181# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2626 a_8837_7983# ts.o_res\[17\] a_8491_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2627 _166_ ts.ts_ctrl.temp_ctr\[5\] a_1775_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2628 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2629 VPWR _058_ a_11573_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2630 VPWR a_4111_4221# a_4279_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2631 VPWR _073_ _094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X2632 a_6515_5108# _221_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2633 a_16170_6895# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X2634 VPWR _065_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X2635 a_6607_17687# ts.ts_ctrl.temp_ctr\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2636 _064_ a_13731_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2637 a_12910_10199# _069_ a_12829_10199# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X2638 net17 a_6559_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2639 a_8907_4182# ts.o_res\[19\] a_8448_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2640 VPWR net4 a_18597_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X2641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2643 VGND a_9287_3829# _154_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2644 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2645 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2646 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2647 a_4515_4399# a_3891_4405# a_4407_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2648 VPWR _059_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2649 net16 a_5423_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2650 a_15308_7369# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2651 a_17051_14997# a_16863_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2652 a_10335_4117# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2653 a_9460_13799# ts.ts_ctrl.temp_ctr\[6\] a_9602_13974# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X2654 uo_out[3] a_8468_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2655 a_7994_13469# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2656 a_6796_17999# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2657 a_6427_16341# _186_ a_6645_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X2658 a_5161_14735# a_4995_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2659 ts.ts_core.dac_vout_ana_ net15 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2660 a_14664_12809# a_15399_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2661 ts.ts_core.dac_vout_ana_ net71 a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2662 VGND net67 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2663 a_10883_4943# _155_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X2664 VGND net69 a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2665 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X2666 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2667 VPWR net68 a_16863_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2668 VPWR _077_ a_12894_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X2669 a_4696_17833# a_3615_17461# a_4349_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2670 VGND a_2751_15253# a_2493_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X2671 VGND ts.ts_ctrl.temp_ctr\[1\] a_10759_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2672 a_14296_4399# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2673 VGND _114_ a_12883_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X2674 a_3299_9269# _163_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X2675 a_1021_14735# a_855_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2676 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2677 VPWR a_12321_12705# _103_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2678 VPWR a_1459_14423# _016_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X2679 a_8468_10357# _055_ a_8856_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2681 a_14475_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2682 VGND _067_ a_14937_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2683 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2684 a_4071_7369# ts.ts_ctrl.temp_ctr\[17\] a_3853_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2685 a_10649_15823# a_10605_16065# a_10483_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2687 a_15123_2197# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2688 VPWR a_3299_12533# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2689 VPWR a_11719_2197# a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X2690 a_13599_6807# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.141 ps=1.33 w=0.42 l=0.15
X2691 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2692 a_7921_2229# a_7755_2229# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2694 VGND net2 a_16771_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X2695 a_12157_9813# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X2696 a_12493_7369# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2697 a_18719_5193# _146_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2698 a_16143_14191# net10 _066_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2699 VPWR a_4588_14709# _177_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2700 VGND ts.ts_ctrl.state\[1\] _112_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2701 a_6244_9117# _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2702 VGND a_7815_13407# a_7749_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2703 VPWR ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_16127_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2704 VGND net70 a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2705 a_17121_4943# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2706 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2708 _182_ ts.ts_ctrl.temp_ctr\[11\] a_7470_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X2709 a_4884_6281# _137_ a_4617_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.165 ps=1.33 w=1 l=0.15
X2710 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2712 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2713 a_9532_18365# a_9095_17973# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2715 a_4341_14557# ts.ts_ctrl.temp_ctr\[8\] a_4259_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X2716 a_15951_2919# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2717 VGND a_7159_16599# _184_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2718 a_13928_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2719 a_10483_15823# a_10037_15823# a_10387_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2720 net55 clknet_2_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2721 a_10200_6031# _008_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2722 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2723 VPWR a_1936_9129# a_2111_9055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2724 VGND a_18937_2932# net7 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2725 a_2397_3855# a_1407_3855# a_2271_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2726 VGND a_14347_3615# a_14281_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2727 VPWR a_3854_3967# a_3781_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2728 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2729 a_11573_7983# _070_ a_11573_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2730 VPWR _094_ a_16407_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X2731 VPWR a_12353_14977# a_12243_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2732 a_1589_10901# a_1371_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2733 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2734 net12 a_18847_16341# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2735 a_14545_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2736 a_11399_1109# ts.ts_core.tempdelay_sync1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2737 VPWR _162_ a_2451_9323# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2738 a_8022_6575# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2739 uo_out[4] a_9340_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X2740 net72 a_18335_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2741 a_9256_11471# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2742 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2743 VGND _201_ a_4956_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X2744 a_5161_14735# a_4995_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2745 a_13832_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2746 a_7109_18241# a_6891_17999# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2747 a_7719_17833# a_7369_17461# a_7624_17821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2748 VPWR a_12547_4007# a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2749 a_16661_11247# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2750 a_5269_15279# _186_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2751 a_11517_9117# ts.ts_ctrl.state\[1\] a_11435_8864# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2752 VPWR ts.ts_ctrl.temp_ctr\[15\] _189_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2753 a_15259_13423# net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2754 VGND net70 a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2755 a_4425_10383# a_4259_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2756 a_12029_17821# a_11985_17429# a_11863_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2757 a_10391_14709# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2758 a_16499_12821# a_16311_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2759 a_8360_15645# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2760 a_15763_4117# a_15575_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2761 a_17673_6895# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2762 a_1021_14735# a_855_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2763 VPWR _140_ a_16589_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.117 ps=1.24 w=1 l=0.15
X2764 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2765 a_18234_10927# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2766 a_9629_13103# _057_ a_9800_13423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2767 a_2493_14197# a_2327_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2768 VGND _047_ a_9256_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2769 a_10313_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2771 a_15959_10633# _068_ _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2772 ts.ts_core.capload\[14\].cap.Y net27 a_6553_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2773 VGND _137_ _201_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.115 ps=1 w=0.65 l=0.15
X2774 _154_ a_9287_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2775 a_16315_13103# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2776 a_4871_17759# a_4696_17833# a_5050_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2777 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2778 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2779 a_6785_6941# a_6741_6549# a_6619_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2780 VGND ts.o_res\[12\] a_9608_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X2781 a_16477_12559# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2782 ts.o_res\[19\] a_7539_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2783 _124_ a_11435_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X2784 a_16960_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2785 ts.ts_ctrl.temp_ctr\[9\] a_2111_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2786 VPWR a_10625_7352# a_10294_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X2787 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2788 VPWR a_17507_4399# a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2789 VGND net70 a_15299_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2790 a_13821_6941# _114_ a_13733_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X2791 VGND _051_ a_11188_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2792 a_16293_13423# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2793 VPWR a_7017_4097# a_6907_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2794 VGND a_13327_9813# _089_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X2795 VGND net68 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2796 _201_ _200_ a_4884_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.35 w=1 l=0.15
X2797 a_15304_7119# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2798 ts.ts_core.dac_vout_ana_ net72 a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2799 net53 clknet_2_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2800 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2801 a_7737_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2802 a_11812_841# a_12547_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2803 a_1467_14735# a_1021_14735# a_1371_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2804 a_13295_11247# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X2805 a_3781_4221# a_3247_3855# a_3686_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2806 VGND _061_ a_16354_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2807 a_1276_9117# _010_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2808 VPWR clknet_2_3__leaf_clk a_11711_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2809 VPWR _061_ a_13643_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X2810 a_14281_10205# a_14011_9839# a_14177_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2811 a_9290_10633# ts.o_res\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X2812 VGND _173_ a_1677_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2813 _143_ _059_ a_13601_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2815 a_12241_13423# ts.ts_ctrl.temp_ctr\[5\] a_11895_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2816 a_4867_12559# a_4351_12559# a_4772_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2817 VPWR a_4687_4917# a_4674_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2818 _050_ net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2819 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2820 VPWR a_12631_2223# a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2821 a_1585_8457# _161_ a_1501_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2822 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2823 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
R30 VPWR ts.ts_core.capload\[14\].cap_27.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2824 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2825 a_9823_13647# ts.ts_ctrl.temp_ctr\[6\] a_9460_13799# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2827 a_17695_15279# a_17507_15279# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X2828 ts.ts_core.dac_vout_ana_ net15 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2829 VPWR ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref a_16955_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2830 VPWR a_4503_8181# a_4490_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2831 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2832 ts.o_res\[16\] a_7263_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2833 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2834 a_14882_7983# _065_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2835 VGND a_9460_13799# _208_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2836 VGND net69 a_14379_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2837 _161_ ts.ts_ctrl.temp_ctr\[2\] a_1858_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X2838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2839 a_6428_6941# _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2840 ts.ts_core.dac_vout_ana_ net47 a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2841 VPWR ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref a_18234_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2842 VPWR a_10147_2767# a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2843 a_1936_12559# a_1021_12559# a_1589_12801# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2844 ts.ts_core.capload\[10\].cap.Y net23 a_7381_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2845 VGND ts.ts_ctrl.temp_ctr\[19\] _200_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2846 a_13845_7369# _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2848 ts.ts_core.dac_vout_ana_ net72 a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2849 VGND a_9771_18236# a_9702_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2851 a_8500_1929# a_9235_1831# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2852 VGND _087_ a_9941_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2853 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14292_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2854 a_12650_12809# _101_ a_12570_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X2855 a_8879_4438# ts.o_res\[0\] a_8807_4438# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2856 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2857 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2858 ts.ts_core.tempdelay_sync1 a_8787_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2859 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2860 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2861 VPWR a_12047_6835# _061_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2862 net69 a_18234_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2863 a_12603_9545# _105_ a_12531_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2864 a_7719_15797# ts.ts_ctrl.temp_ctr\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2865 _201_ _200_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.112 ps=0.995 w=0.65 l=0.15
X2866 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2867 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2868 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_11803_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2869 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2870 a_12267_1135# a_12079_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2871 a_17599_6031# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2872 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2873 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2874 a_9503_9295# _088_ a_9681_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2875 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2876 ts.ts_core.dac_vout_ana_ net15 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2877 ts.ts_core.dac_vout_ana_ net14 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2878 a_18774_3311# a_18597_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X2879 a_17673_15599# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2880 a_10313_2767# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2881 VGND a_13231_12247# _081_ VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2882 a_2375_12247# _164_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X2883 VGND a_10275_4399# a_10443_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2884 a_9869_14977# a_9651_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2885 a_16129_4399# ts.ts_ctrl.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2886 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2887 a_6839_853# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2888 VPWR clknet_2_3__leaf_clk a_6559_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2889 a_7117_14735# _177_ a_7045_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2890 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2891 VGND a_8175_3285# ts.o_res\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2892 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2893 a_11601_4943# ts.ts_ctrl.state\[1\] a_11517_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X2894 a_12679_10071# a_12952_10071# a_12910_10199# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2895 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2896 _198_ a_4075_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2897 VPWR a_13326_5719# _146_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X2898 _171_ a_2787_10205# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X2899 a_4135_11445# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2900 VPWR _050_ a_11359_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2901 a_16775_7663# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2902 VGND _120_ a_11236_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
X2903 a_8695_3553# clknet_2_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2905 a_11808_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2906 a_16499_12821# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2907 VGND net17 a_6785_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2908 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2909 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2910 a_10478_16911# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2911 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2912 a_1276_12559# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2913 VPWR a_6883_14887# _186_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2914 a_8679_3029# a_8491_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2915 a_12547_4007# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2916 a_12679_10071# a_12952_10071# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2917 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2918 VPWR _065_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2919 VPWR a_5432_12559# a_5607_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2920 VGND net68 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2922 _023_ _194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2923 VGND _166_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2924 a_13901_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2925 VPWR _156_ a_11255_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2926 VGND net69 a_17507_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2927 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2928 VPWR a_5043_13322# _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2929 VPWR a_14295_2919# a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2930 a_9287_3829# _153_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2931 a_18836_12711# net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.321 ps=1.68 w=0.42 l=0.15
X2932 a_4073_14985# ts.ts_ctrl.temp_ctr\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2933 a_14471_8207# _059_ _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2934 a_9275_6358# ts.o_res\[1\] a_8816_6183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2935 VGND a_7079_7967# a_7013_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2936 a_14195_9545# _133_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2937 VPWR _084_ a_11877_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2938 VGND _211_ a_11753_16150# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X2939 a_17121_14511# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2940 _094_ a_15535_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2941 VPWR a_9227_2223# a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2942 a_1633_9117# a_1589_8725# a_1467_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2943 a_8455_15657# a_7939_15285# a_8360_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2945 ts.ts_core.dac_vout_ana_ net15 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2946 VGND _120_ a_11159_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2947 a_3571_16586# _180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2948 ts.ts_core.dac_vout_ana_ net15 a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X2949 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2950 a_7221_7093# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2951 VPWR ts.ts_ctrl.temp_ctr\[13\] a_6998_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X2952 a_16591_1135# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2953 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2954 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2955 a_4393_17821# a_4349_17429# a_4227_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2956 a_17029_14735# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2957 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X2958 a_14475_5205# a_14287_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2960 _092_ a_9503_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2961 VPWR clknet_2_2__leaf_clk a_2879_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2962 VGND a_2439_4123# a_2397_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2963 VGND a_11851_12247# _116_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2964 ts.ts_core.dac_vout_ana_ net71 a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2965 VPWR a_12777_6005# _144_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2966 _084_ a_12603_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2967 a_3111_6794# _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2968 VGND a_4503_8181# a_4437_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2969 a_6723_15279# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2970 a_13845_7369# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2971 _029_ a_5455_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2972 a_7221_7093# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2973 a_10239_9295# _088_ a_10417_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2974 a_3413_15823# a_3247_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2975 VGND ts.ts_core.dac.vdac_single.en_pupd a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2976 VPWR ts.ts_ctrl.temp_ctr\[12\] a_6607_17687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2977 VGND clknet_2_0__leaf_clk a_3891_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2978 _130_ a_9214_10159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2979 a_2537_12381# _164_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X2980 _061_ a_12047_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2981 a_13923_1135# a_13735_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X2982 a_13365_12381# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.103 ps=1 w=0.42 l=0.15
X2983 VPWR a_14584_8751# uio_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2984 a_14526_14165# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2985 ts.ts_core.tempdelay_async ts.ts_core.dcdel_out_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2986 a_4866_4943# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2987 a_11875_17455# a_11251_17461# a_11767_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2988 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2989 VGND net69 a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2990 a_13599_6807# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X2991 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2992 a_1276_9117# _010_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2993 VPWR a_4165_5185# a_4055_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2994 VPWR a_14379_6575# a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X2995 VGND clknet_2_2__leaf_clk a_4995_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2996 a_12079_8457# _124_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2997 a_16569_10383# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2998 a_17143_8469# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2999 VGND _125_ a_12851_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3000 ts.o_res\[6\] a_10391_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3001 VPWR clk a_7286_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3002 a_17935_13363# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3003 a_7759_1135# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3004 a_7456_17999# a_6375_17999# a_7109_18241# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3005 _093_ a_10977_9955# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3006 a_5271_13216# ts.ts_ctrl.temp_ctr\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3007 a_4365_9111# _192_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.13 ps=1.11 w=0.42 l=0.15
X3008 a_9770_10633# ts.o_res\[16\] a_9687_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3009 a_14660_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3010 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _061_ a_16793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3012 net67 a_17332_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3013 _006_ a_16298_4719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X3014 a_7442_4765# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3016 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3017 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3018 VPWR a_16587_7663# a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3019 a_9747_14735# a_9301_14735# a_9651_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3020 a_6331_12234# _209_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3022 _076_ a_9770_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X3023 a_6181_591# net28 ts.ts_core.capload\[15\].cap.Y VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3024 a_13834_8207# net7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.12 ps=1.04 w=0.65 l=0.15
X3025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3026 a_15649_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3027 a_13560_841# a_14295_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3028 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_17783_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3029 ts.ts_core.dac_vout_ana_ net15 a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3030 VGND clknet_2_1__leaf_clk a_6283_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3031 VGND a_7355_15583# a_7289_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3032 VGND a_8448_4007# _222_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3033 VGND _135_ a_14195_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3035 a_6239_8534# ts.o_res\[3\] a_5780_8359# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X3036 a_15216_3017# a_15951_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X3037 VGND net69 a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3038 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3039 VPWR ts.ts_ctrl.temp_ctr\[10\] a_5271_13216# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3040 VPWR ts.ts_ctrl.temp_ctr\[17\] _196_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3041 VPWR a_18755_3829# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3042 VPWR _098_ a_13741_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3043 VGND net69 a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3044 a_9971_743# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3045 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3046 a_17603_9839# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3047 _148_ a_17753_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3048 VPWR a_16495_12015# a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3049 a_17121_7119# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3050 _177_ a_4588_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3051 a_11626_17238# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3052 a_9232_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3053 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X3054 a_1367_10357# _165_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X3055 _019_ _183_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3056 VGND a_6209_8181# a_6143_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3057 a_11679_6183# _062_ a_11853_6059# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3058 a_6607_17687# ts.ts_ctrl.temp_ctr\[11\] a_6841_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3059 a_8679_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3060 a_3701_8751# _193_ a_3617_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3061 VGND a_11760_14423# _212_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3062 a_11969_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3063 a_13556_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3064 a_5085_5487# _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X3065 a_10141_6575# _112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X3066 _065_ _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3067 a_9232_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3068 a_14471_13423# net11 _059_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3069 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3070 VPWR a_15031_4373# a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3071 net68 a_13611_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3072 a_17753_9545# net3 a_17599_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X3073 a_14353_10205# _068_ a_14281_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3074 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3075 VGND _050_ _122_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3076 a_13928_5487# a_14663_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3077 a_1479_7485# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3078 VGND a_2111_14709# ts.ts_ctrl.temp_ctr\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3079 VPWR ts.ts_ctrl.temp_ctr\[2\] a_2755_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3080 uo_out[2] a_11272_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3081 VGND a_11478_4373# a_11119_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3082 VPWR a_8632_16599# _214_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3083 VPWR _139_ a_11467_5825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3084 _073_ a_16640_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3085 a_11991_1941# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3086 VPWR a_8836_10901# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3088 a_18243_7663# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3089 a_15952_9545# a_16687_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3090 a_4513_13621# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3091 VGND a_5043_13322# _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3092 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3093 a_17143_5205# a_16955_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3094 a_11808_4943# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3095 VPWR _177_ a_7387_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X3096 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3098 ts.ts_core.dac_vout_ana_ net14 a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3099 VPWR net34 ts.ts_core.capload\[6\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3100 a_4682_15823# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3101 a_10980_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3102 a_4195_4221# a_3413_3855# a_4111_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3103 VPWR clknet_2_2__leaf_clk a_4995_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3104 a_9582_12335# ts.o_res\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X3105 a_9615_18141# clknet_2_3__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3106 a_2701_13897# _173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3107 ts.o_res\[11\] a_10299_16885# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3108 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3109 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd a_12997_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X3110 a_9224_10927# _049_ a_8836_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X3111 VGND net13 a_15259_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3112 _189_ ts.ts_ctrl.temp_ctr\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3113 a_13463_5807# net4 a_13326_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3114 VGND a_4956_5461# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X3115 VPWR _069_ a_9687_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X3116 VGND net8 _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3117 VPWR a_16311_12559# a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3118 VPWR a_10147_1679# a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3119 a_16293_13423# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3120 a_12691_7663# _122_ a_12597_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X3121 a_9655_16911# a_9209_16911# a_9559_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3122 a_14545_6895# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3124 a_9393_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3125 a_3299_12533# _167_ a_3517_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X3126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3127 a_9800_13423# net8 a_9629_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X3128 VPWR clknet_2_1__leaf_clk a_6283_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3129 a_13595_12336# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3130 VPWR clknet_2_2__leaf_clk a_2327_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3131 VPWR a_13059_4703# ts.ts_ctrl.state\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3132 VPWR a_16403_1135# a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3133 a_16477_12559# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3134 a_11484_17063# ts.ts_ctrl.temp_ctr\[13\] a_11626_17238# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X3135 _059_ net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3136 a_4625_4373# a_4407_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3137 VPWR a_4871_17759# ts.ts_ctrl.temp_ctr\[11\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3138 a_17051_3029# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3139 a_9679_9955# _132_ a_9597_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3140 a_4617_6281# _194_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3141 a_7066_8751# a_5989_8757# a_6904_9129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3142 a_16591_10645# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3143 a_15259_13423# net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3144 a_9608_11471# _051_ a_9340_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3145 a_8415_13103# net9 _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3146 VGND a_4503_15797# a_4437_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3147 _096_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_18243_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3148 a_4713_16911# net63 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3149 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3150 VGND a_10443_4373# a_10401_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3151 VGND net70 a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3152 a_11188_11471# ts.o_res\[10\] a_11272_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3153 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3154 a_14935_1941# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3155 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_10147_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3156 _053_ a_7775_8534# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3157 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3158 a_13556_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3159 VPWR a_17507_6575# a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3160 a_19057_3311# a_18880_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3161 VPWR a_5893_17687# net63 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3162 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3163 a_9770_9071# ts.ts_ctrl.temp_ctr\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X3164 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3165 a_12243_15101# a_11619_14735# a_12135_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3166 VPWR a_6607_17687# _183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3167 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3168 a_6883_14887# ts.ts_ctrl.state\[2\] a_7117_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3169 a_15308_7369# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3170 ts.ts_core.dac_vout_ana_ net14 a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3171 a_14567_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3172 a_5269_15279# net58 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3173 a_10335_4117# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3175 ts.ts_core.dac_vout_ana_ net15 a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3176 a_11035_6005# a_10860_6031# a_11214_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3177 a_17121_14511# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3178 VPWR a_16955_14191# a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3179 VGND _061_ a_16170_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3180 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3181 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3182 VGND net17 a_13869_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3183 a_11606_7119# _058_ a_11520_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X3184 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3185 a_4239_17455# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3186 a_18969_5487# _148_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3187 a_2111_7093# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3188 VGND a_5780_8359# _205_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3189 VPWR a_17507_8751# a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3190 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3192 a_9629_13103# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X3193 a_15031_4373# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3194 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
D0 VGND ui_in[2] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X3195 VPWR a_7571_1135# a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3196 VPWR a_6516_11159# _209_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3197 a_7203_12015# net21 a_7285_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3198 ts.ts_core.dac_vout_ana_ net47 a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3199 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3200 VPWR _069_ a_11435_8864# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3201 VGND _147_ a_15943_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3202 a_2929_9089# ts.ts_ctrl.temp_ctr\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X3203 a_14475_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3204 a_6839_853# a_6651_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3206 VPWR ts.ts_ctrl.state\[2\] a_4071_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3207 a_9577_4405# a_9411_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3208 VPWR a_13503_10145# a_13327_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X3209 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3210 a_8468_10357# net8 a_8938_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3211 a_17143_14191# a_16955_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X3212 a_16109_6031# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3213 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3214 VPWR _075_ a_7929_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3215 a_8362_2197# a_8194_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3217 a_5694_10383# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3218 a_8235_8790# ts.o_res\[19\] a_8163_8790# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3219 VPWR a_6059_6005# _137_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3220 a_14687_13693# net13 a_14583_13693# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X3221 VGND _154_ a_9100_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X3222 VPWR a_15943_6031# a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3223 _170_ _164_ a_2778_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X3224 VPWR a_17415_9839# a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3225 a_9236_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3226 uio_out[6] a_12127_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3227 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3228 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3229 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3230 a_17332_3829# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3231 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3232 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3233 a_8879_4438# ts.ts_ctrl.temp_ctr\[0\] a_8879_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3234 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3235 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3236 VGND _127_ a_10975_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X3237 a_12819_2223# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3238 a_16109_6031# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3239 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3240 VGND _141_ a_18821_6059# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3241 VPWR a_7252_12711# _207_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3242 VPWR _068_ a_13086_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X3243 a_14085_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3244 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3245 VPWR _114_ _174_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3246 a_12547_5095# net68 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3247 a_11975_5461# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3248 a_7203_12015# net21 a_7285_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3249 VGND net20 a_4393_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3250 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3252 a_17143_5205# a_16955_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X3253 a_10313_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3254 net65 a_15571_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3255 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3256 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3257 a_14296_4399# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3258 a_9195_15583# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3259 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref _150_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3260 a_1936_14735# a_855_14735# a_1589_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3261 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3262 a_16640_14165# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3263 ts.ts_core.capload\[14\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3264 a_1589_10901# a_1371_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3266 a_11573_7983# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3267 VGND a_5515_10357# a_5449_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3268 a_6601_11471# a_6557_11713# a_6435_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3269 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3270 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3271 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
R31 VPWR ts.ts_core.capload\[10\].cap_23.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3272 a_6817_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3273 a_10965_5193# _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X3274 VPWR a_10147_1679# a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3275 a_7737_1455# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3276 a_17695_4399# a_17507_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3277 a_9415_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3278 VPWR _211_ a_11753_16150# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X3279 a_16315_853# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3280 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_13183_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3281 VPWR a_14717_9545# uio_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3282 VGND net69 a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3283 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3284 a_13556_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3285 a_14913_1679# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3286 a_16569_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3287 a_7079_7967# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3288 a_17673_6895# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3289 a_10138_10927# ts.o_res\[7\] a_10055_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3290 a_13607_3689# a_13091_3317# a_13512_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3291 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3292 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3293 a_14567_12015# a_14379_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3294 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3295 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3296 a_12445_15253# a_12227_15657# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3297 ts.ts_ctrl.temp_ctr\[16\] a_4503_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3298 ts.ts_ctrl.temp_ctr\[10\] a_4503_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3299 a_8853_5865# a_7663_5493# a_8744_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3300 VGND a_8468_10357# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3301 VPWR ts.ts_ctrl.state\[2\] a_15229_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3302 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3303 a_9415_1135# a_9227_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3304 VPWR net59 a_4684_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X3305 _169_ _164_ a_2873_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3306 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.capload\[8\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3307 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3308 a_15763_4117# a_15575_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3310 a_17029_1679# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3311 a_1371_11305# a_1021_10933# a_1276_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3312 VGND net19 a_7153_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3313 a_18755_3829# _142_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X3314 VGND a_13059_4703# ts.ts_ctrl.state\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3315 VPWR _200_ a_5085_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3316 a_10239_13897# _082_ a_10321_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3317 VPWR a_6557_8725# a_6447_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3318 VPWR _067_ a_13231_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X3319 _130_ a_9214_10159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X3320 a_5607_12533# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3321 VGND _187_ a_6153_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.266 pd=2.12 as=0.091 ps=0.93 w=0.65 l=0.15
X3322 _012_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3323 VGND a_9615_18141# a_9576_18267# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3324 a_10313_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3325 a_9777_17153# a_9559_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3326 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3327 VPWR _074_ a_14063_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X3328 a_16683_12015# a_16495_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
R32 uio_oe[4] VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3329 a_9850_4399# a_9411_4405# a_9765_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3330 a_2951_14191# a_2327_14197# a_2843_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3331 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3332 a_17051_14997# a_16863_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
R33 net37 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3333 VPWR a_16863_1679# a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3334 ts.ts_core.capload\[10\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3335 VPWR a_15123_2197# a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3336 a_9098_5853# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3337 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3338 a_13836_11721# a_14571_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3339 a_1371_12559# a_855_12559# a_1276_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3340 a_15304_7119# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3341 ts.ts_core.dac_vout_ana_ net72 a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3342 a_7737_1455# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3343 _110_ _109_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3344 VGND _117_ a_11343_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3345 VPWR a_5179_16367# _138_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3346 VGND a_9287_3829# _154_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3347 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3348 net20 a_4680_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3349 a_9277_8534# ts.o_res\[1\] a_9063_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X3350 a_14295_743# net67 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3351 a_13101_7369# _111_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3353 VPWR a_8619_2223# a_8787_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3355 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3357 a_10055_10927# _088_ a_10138_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X3358 VPWR _168_ a_2695_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X3359 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3360 a_13845_7369# _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3361 ts.ts_core.dac_vout_ana_ net15 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3362 VPWR clknet_2_0__leaf_clk a_3431_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3363 a_10625_7352# ts.ts_ctrl.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X3364 _104_ a_11435_8864# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3365 VPWR clknet_2_2__leaf_clk a_855_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3366 VPWR clknet_2_2__leaf_clk a_3247_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3367 VGND ts.ts_ctrl.temp_ctr\[8\] a_3247_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3368 ts.ts_core.dac_vout_ana_ net14 a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3369 VGND net67 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3370 a_12884_4777# a_11969_4405# a_12537_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3371 VPWR _067_ a_14011_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3373 a_11159_13103# _081_ a_11337_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3374 a_13059_4703# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3375 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3376 ts.o_res\[5\] a_7815_13407# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3377 VPWR a_10441_5785# a_10471_5526# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3378 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3379 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3380 a_8745_7119# ts.o_res\[18\] a_8399_7369# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3381 a_18325_9545# _141_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3382 VPWR a_10011_3530# _027_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3383 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3384 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3385 VPWR a_10147_2767# a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3386 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3387 a_16661_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3388 ts.ts_core.dac_vout_ana_ net72 a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3389 VGND net70 a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3390 net67 a_17332_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3391 _155_ a_10523_3427# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X3392 _122_ _059_ a_12631_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3393 a_3854_3967# a_3686_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3394 net4 a_18278_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3396 VPWR a_11484_17063# _216_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3397 VGND a_6629_15975# net58 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3398 a_8500_1929# a_9235_1831# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3399 VGND net69 a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3400 a_5147_4703# a_4972_4777# a_5326_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3401 a_16499_12821# a_16311_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X3402 a_13755_13423# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X3403 a_7337_13469# a_7293_13077# a_7171_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3404 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _065_ a_14882_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3405 a_16771_10159# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3407 _015_ _174_ a_2701_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3408 a_7180_15657# a_6265_15285# a_6833_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3409 a_5416_14735# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3410 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15575_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3411 a_13546_10535# a_14015_10357# a_13959_10429# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X3412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3413 a_17121_4943# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3414 VPWR a_2111_7093# a_2098_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3415 a_10689_12809# ts.o_res\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3416 a_4975_12925# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3417 a_10037_15823# a_9871_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3418 ts.o_res\[4\] a_5515_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3419 a_10830_10633# _070_ a_10516_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X3420 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3421 net9 a_18671_14451# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3422 a_9976_4777# a_9577_4405# a_9850_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3423 a_3613_10901# a_3395_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3424 VGND net16 a_6601_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3425 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3426 a_3671_12393# a_3321_12021# a_3576_12381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3427 ts.ts_core.dac_vout_ana_ net14 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3428 ts.ts_core.dac_vout_ana_ net15 a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X3429 a_8933_4943# a_8767_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3430 VGND _091_ a_9503_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3431 a_7079_7967# a_6904_8041# a_7258_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3432 a_16569_10383# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3433 a_7180_15657# a_6099_15285# a_6833_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3434 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3435 VGND clknet_2_3__leaf_clk a_9871_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3436 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3437 a_16683_12015# a_16495_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3438 ts.ts_core.dac_vout_ana_ net14 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3439 a_13551_6031# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3440 a_7681_12533# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3441 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3442 a_15741_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3443 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9227_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3444 a_9209_16911# a_9043_16911# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3446 a_11599_3311# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3447 a_13715_3311# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3448 VGND a_12189_14489# a_12123_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3449 VPWR ts.ts_ctrl.temp_ctr\[13\] a_6427_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X3450 a_9957_3855# _062_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3451 ts.o_res\[15\] a_9195_15583# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3453 VPWR _055_ a_8938_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X3454 uio_out[7] a_14717_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3455 VGND a_17191_11445# _074_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3456 a_17029_1679# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3457 VPWR _067_ a_13445_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X3458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3459 a_7681_12533# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X3460 ts.o_res\[18\] a_7263_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3461 a_16775_7663# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3462 VPWR ts.o_res\[8\] a_9687_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X3463 _123_ a_8399_7369# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3464 VGND a_1551_6807# _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3465 VPWR _147_ a_15943_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3466 VGND a_2271_4221# a_2439_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3467 VGND net69 a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3468 a_8284_17833# a_7203_17461# a_7937_17429# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3469 _182_ ts.ts_ctrl.temp_ctr\[12\] a_7387_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3470 a_18763_9447# _099_ a_18937_9323# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3471 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3472 _215_ a_9339_18582# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3473 ts.ts_core.tempdelay_sync1 a_8787_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3474 a_13963_6896# _095_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3475 VPWR a_1936_11305# a_2111_11231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3476 VGND a_6884_5095# _221_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X3477 VPWR a_9848_4943# a_10023_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3478 a_2098_8751# a_1021_8757# a_1936_9129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3479 a_8907_9622# ts.o_res\[16\] a_8448_9447# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X3480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3481 ts.ts_core.capload\[7\].cap.Y net35 a_6921_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3482 a_16687_9447# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3483 a_14986_9849# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X3484 _023_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3485 a_13901_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3486 a_14347_3615# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3487 a_15465_13647# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3488 VGND clknet_0_clk a_4513_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3489 VPWR ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_13919_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3490 VPWR a_14295_2919# a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3491 a_11895_13103# _082_ a_11977_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3492 VPWR a_8836_10901# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3493 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
R34 uio_oe[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3494 a_8573_7663# ts.o_res\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3495 a_14418_9071# _100_ a_14584_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3496 a_16293_13423# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3497 a_17581_10159# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3498 _120_ a_10975_8864# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3499 VGND _062_ a_12275_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X3500 a_7847_12015# net21 a_7929_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3502 _004_ a_11056_5193# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3503 VGND net55 a_9411_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3504 a_15308_8457# net47 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3505 a_16293_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3506 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3507 VPWR a_9227_2223# a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3508 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3509 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3510 a_10154_15318# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3511 VPWR res1_n a_3177_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3512 a_9283_4943# a_8933_4943# a_9188_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3513 a_3413_3311# a_3177_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X3514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3515 VGND _137_ a_5232_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X3516 a_11606_7119# net7 a_11437_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X3517 _121_ a_11159_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X3518 a_16591_1135# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3519 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3520 VPWR net67 a_15943_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3521 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3522 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3523 a_14374_13799# a_14733_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3524 VPWR clknet_2_0__leaf_clk a_5823_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3525 VPWR _115_ a_12329_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3526 a_14475_5205# a_14287_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3527 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3528 a_4236_12393# a_3155_12021# a_3889_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3529 a_3663_15511# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3530 VPWR a_12547_5095# a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3531 ts.ts_ctrl.temp_ctr\[11\] a_4871_17759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3532 a_12227_15657# a_11711_15285# a_12132_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3533 a_15159_11248# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3534 ts.ts_core.dac_vout_ana_ net71 a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3535 VPWR net12 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3537 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X3538 a_14063_10901# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X3539 _068_ a_13603_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3540 VPWR a_10147_2767# a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3541 _047_ net9 a_8415_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3542 a_13845_7369# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3543 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3544 a_6904_9129# a_5989_8757# a_6557_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3545 a_17783_5487# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3546 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd _061_ a_17034_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.175 ps=1.35 w=1 l=0.15
X3547 a_3571_16586# _180_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3548 a_16964_13897# a_17699_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3549 a_12132_15645# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3550 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10335_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X3551 net14 a_17783_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3552 VPWR ts.ts_ctrl.temp_ctr\[2\] a_11610_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3553 _196_ _194_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3554 VGND a_10011_3530# _027_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3555 a_15304_7119# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3556 VPWR _139_ a_18763_7271# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3557 a_11429_6941# a_11159_6575# a_11339_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3558 a_11425_12809# _118_ a_11343_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X3559 VGND a_7079_11445# a_7013_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3560 a_12809_14735# a_11619_14735# a_12700_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3562 VPWR a_14584_8751# uio_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3563 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3564 a_13546_13335# a_13905_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3565 a_7802_13103# a_6725_13109# a_7640_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3567 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3568 VGND net18 a_6601_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3570 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3571 a_3111_6794# _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3572 a_4157_6031# ts.ts_ctrl.state\[2\] a_4075_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3573 a_5381_11225# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X3574 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3575 a_9236_841# a_9971_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X3576 a_4963_12559# a_4517_12559# a_4867_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3577 a_17143_14191# a_16955_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3578 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3579 VPWR a_4329_13335# net62 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3580 a_16315_2223# a_16127_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3581 VGND clknet_2_0__leaf_clk a_6007_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3582 a_6999_18365# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3583 ts.ts_core.dac_vout_ana_ net72 a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3584 VGND net67 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3585 a_16591_10645# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3586 VPWR a_14295_743# a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3587 VPWR a_12047_6835# _061_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3588 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3589 VPWR a_14063_10901# _077_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X3590 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3591 a_7759_1135# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3594 a_6791_3530# _222_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3595 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3596 a_7251_7446# ts.o_res\[2\] a_6792_7271# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X3597 VGND _071_ a_10493_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3598 ts.ts_ctrl.temp_ctr\[0\] a_10023_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3599 _168_ a_2695_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3600 VGND a_2111_7093# a_2045_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3601 a_14453_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3602 ts.o_res\[10\] a_12967_15583# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3603 uo_out[5] a_9524_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3604 a_1021_10933# a_855_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3605 VPWR a_16863_2767# a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3606 a_3671_12393# a_3155_12021# a_3576_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3607 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3608 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3609 a_3045_10933# a_2879_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3611 a_10012_15511# ts.ts_ctrl.temp_ctr\[14\] a_10154_15318# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X3612 VPWR a_4236_12393# a_4411_12319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3614 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3615 a_16793_8751# _061_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3616 a_17121_14511# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3617 a_8679_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3618 VPWR a_16955_14191# a_17143_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3619 VGND a_7221_7093# a_7155_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3620 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3621 VPWR _191_ a_5871_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3622 VPWR _065_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3623 a_6607_17687# _177_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3624 a_9391_5309# a_8767_4943# a_9283_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3625 ts.ts_core.capload\[4\].cap.Y net32 a_7105_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3626 VPWR a_11975_5461# net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3627 a_12686_17821# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3628 a_11991_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3629 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3630 VPWR _177_ a_6067_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3631 VPWR net13 a_13905_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X3632 a_16170_6895# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3633 a_4517_12559# a_4351_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3634 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3635 VPWR net10 a_14526_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X3636 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12079_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3637 VPWR _205_ a_5363_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3638 a_16499_12821# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3639 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3640 _211_ a_7815_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3641 a_12219_14230# ts.o_res\[9\] a_11760_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X3642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3643 _094_ _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X3644 _119_ a_11343_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X3645 a_18848_13621# uio_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3646 a_8679_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3647 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3648 a_17143_8469# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3649 a_18109_10548# _152_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3650 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3651 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3652 VPWR a_15031_4373# a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3654 VGND a_12321_12705# _103_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X3655 VGND ts.ts_core.dac_vout_ana_ a_13643_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3656 a_7631_17973# a_7456_17999# a_7810_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3657 a_8496_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3658 a_6904_8041# a_5989_7669# a_6557_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3659 VPWR a_1589_8725# a_1479_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3660 VGND a_9095_17973# ts.o_res\[12\] VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3661 VPWR a_16863_14735# a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3662 ts.ts_core.capload\[6\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3663 a_13928_5487# a_14663_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3664 a_3061_14165# a_2843_14569# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3665 a_3947_4943# a_3597_4943# a_3852_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3666 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3667 VPWR a_8877_3829# a_8907_4182# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3668 a_6631_6575# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3669 VPWR a_14287_6031# a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3670 a_8217_10927# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3671 ts.ts_core.dac_vout_ana_ net14 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3672 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3673 a_11808_3855# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3674 VPWR a_13611_4917# net68 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3675 a_18243_7663# _095_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3676 VPWR a_9227_2223# a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3677 a_3763_8207# a_3413_8207# a_3668_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3678 VGND a_12507_17759# a_12441_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3679 a_14453_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3680 a_10387_15823# a_10037_15823# a_10292_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3681 VGND a_10294_7093# _159_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3682 VGND net12 a_14733_13799# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X3683 a_16569_10383# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3684 a_3063_10205# _162_ a_2957_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3688 VPWR a_2111_11231# ts.ts_ctrl.temp_ctr\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3689 a_3854_3967# a_3686_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3690 a_17121_7119# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3691 VPWR a_14379_12015# a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3692 a_17051_14997# a_16863_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3693 VPWR _061_ a_13769_6296# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.129 ps=1.18 w=0.42 l=0.15
X3694 a_14015_13077# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X3695 VGND clknet_2_0__leaf_clk net52 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3697 uo_out[3] a_8468_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3698 a_13836_11721# a_14571_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3700 _194_ a_4126_8983# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3701 a_11969_2767# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3703 _190_ _189_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X3704 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3705 VPWR a_14331_12533# a_13967_12711# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X3706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3707 VPWR a_16403_1135# a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3708 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3709 a_13901_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3710 VPWR a_14374_13799# _071_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X3711 a_4362_5603# _199_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X3712 a_4775_10383# a_4425_10383# a_4680_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3713 a_12894_10927# _078_ a_12591_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3714 VPWR a_16495_12015# a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3715 a_12056_3689# a_11141_3317# a_11709_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3716 a_14172_3689# a_13257_3317# a_13825_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3717 a_6059_6005# _136_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X3718 net8 a_8399_18543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3719 VPWR a_11272_11471# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3720 a_3713_6941# _195_ a_3641_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3721 a_12809_11247# ts.ts_core.o_tempdelay a_12591_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3722 a_2493_14197# a_2327_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3723 VPWR a_14347_3615# a_14334_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3724 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3725 net16 a_5423_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3726 _096_ _095_ a_18243_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3727 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3728 VPWR a_14379_6575# a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3729 a_8551_15657# a_8105_15285# a_8455_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3730 a_11808_3855# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3731 a_15952_9545# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3733 VPWR a_17507_6575# a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3734 VGND net68 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3735 a_10080_10383# _072_ a_9960_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X3736 VPWR a_18937_11636# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3737 a_16143_14191# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3738 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3739 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3740 a_8500_1929# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3741 a_12829_10199# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X3742 VPWR _075_ a_8573_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3743 a_9667_17277# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3744 VGND net70 a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3745 VGND a_4683_13077# a_4425_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X3746 a_16315_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3747 a_6791_3530# _222_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3748 a_4446_9111# _172_ a_4365_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X3749 VGND clknet_2_3__leaf_clk a_11711_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3750 net67 a_17332_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3751 VPWR a_17507_8751# a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3752 VGND _071_ a_10677_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3753 VGND a_5140_15253# _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X3754 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16587_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3755 a_3871_8573# a_3247_8207# a_3763_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3757 a_7263_6879# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3758 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3759 _161_ ts.ts_ctrl.temp_ctr\[3\] a_1775_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3760 ts.ts_core.dac_vout_ana_ net47 a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3761 a_14331_12533# net12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3762 a_6339_9129# a_5823_8757# a_6244_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3763 VGND clknet_2_1__leaf_clk net54 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3764 a_13183_7663# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3765 VPWR clknet_2_2__leaf_clk a_4259_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3766 a_12954_15279# a_11877_15285# a_12792_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3767 a_3425_5865# a_2235_5493# a_3316_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3768 a_6173_6581# a_6007_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3769 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3770 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3771 a_8397_5461# a_8179_5865# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3772 VGND net69 a_16403_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3773 ts.o_res\[1\] a_8919_5791# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3774 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3775 a_12441_17833# a_11251_17461# a_12332_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3776 a_10605_16065# a_10387_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3777 a_11589_9117# _089_ a_11517_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3778 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3779 a_14857_14342# net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X3780 VPWR net9 a_7981_8790# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X3781 VPWR a_12596_5461# _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3782 a_4713_8751# ts.ts_ctrl.temp_ctr\[16\] _193_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3783 a_11131_9955# _086_ a_11059_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3784 VPWR a_15943_6031# a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3785 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3786 VPWR a_17415_9839# a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X3787 ts.ts_core.dac_vout_ana_ net15 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3788 a_16753_7983# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3789 _069_ _068_ a_15959_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3791 a_10239_13897# _082_ a_10321_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3792 a_8459_17759# a_8284_17833# a_8638_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3793 a_6999_18365# a_6375_17999# a_6891_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3794 VPWR ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14287_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3795 a_10124_16911# a_9043_16911# a_9777_17153# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3796 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3797 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3798 net9 a_18671_14451# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X3799 VGND a_13326_5719# _146_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3800 a_4071_7369# _194_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3801 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3802 a_6076_14735# a_4995_14735# a_5729_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3803 VPWR a_6884_6183# _220_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X3804 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3805 a_14085_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3806 _065_ _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3807 net15 a_11975_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3808 a_5340_10383# a_4259_10383# a_4993_10625# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3809 VGND net16 a_6785_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3810 ts.ts_core.capload\[1\].cap.Y net29 a_6829_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3811 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3812 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3813 a_11808_4943# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3814 a_12591_6895# _112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3815 uo_out[1] a_11456_11247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X3816 a_11325_13103# ts.ts_ctrl.temp_ctr\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3817 a_1479_15101# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3818 VGND net67 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X3819 VPWR net54 a_7755_2229# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3820 a_6799_3855# a_6283_3855# a_6704_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3821 a_14296_4399# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3822 VGND _079_ a_10686_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X3823 ts.ts_core.dac_vout_ana_ net14 a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3824 a_12415_4777# a_11969_4405# a_12319_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3825 _164_ a_3299_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3826 a_15959_10633# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3827 a_16315_13103# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3828 VGND a_3663_15511# _180_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X3829 a_9869_14977# a_9651_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3830 VGND _154_ a_10331_3671# VGND sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X3831 a_7026_6031# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3832 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3833 a_12079_8457# _119_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3834 ts.ts_ctrl.temp_ctr\[9\] a_2111_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3835 uio_out[4] a_11207_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3836 a_17121_7119# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3837 a_6173_9295# a_6007_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3838 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3839 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3840 a_15952_9545# a_16687_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X3841 VGND a_6515_10058# _043_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3842 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3843 VGND net19 a_9333_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X3844 VPWR a_15483_11471# a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3846 a_5050_17821# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3847 a_8938_10633# net8 a_8468_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3848 VPWR a_9889_13621# a_9919_13974# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3849 VPWR a_14717_9545# uio_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3850 a_15465_13647# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3851 a_13556_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3852 a_14913_1679# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3853 a_17029_1679# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3854 _066_ net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3855 a_3657_11293# a_3613_10901# a_3491_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3856 ts.ts_ctrl.state\[0\] a_12231_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3857 ts.ts_ctrl.state\[2\] a_14347_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3858 a_11991_1941# a_11803_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3859 VGND a_11456_11247# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3860 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3861 _080_ a_10686_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X3862 VPWR a_3479_6807# _197_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3863 a_14937_9955# a_14986_9849# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3864 a_2111_12533# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3865 VPWR a_12493_7369# a_12127_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3866 VGND net6 a_14882_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3867 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3868 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3869 a_4219_5461# a_4362_5603# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X3870 a_8744_5865# a_7663_5493# a_8397_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3871 a_15763_4117# a_15575_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3873 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3874 VPWR a_10124_16911# a_10299_16885# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3875 a_10018_4373# a_9850_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3876 a_6339_8041# a_5823_7669# a_6244_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3877 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3878 a_13836_11721# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3879 a_17029_1679# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3880 a_13560_841# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3881 a_14085_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3882 VGND ts.ts_core.dcdel_capnode_ana_ ts.ts_core.dcdel_out_n VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3883 a_2451_9323# _159_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3884 VPWR a_7088_4777# a_7263_4703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3885 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10147_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3886 a_11808_4943# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3887 VGND _158_ _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3888 a_12603_12247# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X3889 a_4126_8983# _192_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.151 ps=1.35 w=0.42 l=0.15
X3890 a_16683_10927# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3891 a_5043_11636# _206_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3892 VGND net70 a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3893 VPWR a_5340_10383# a_5515_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3894 _181_ _137_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3895 a_4517_12559# a_4351_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3896 a_10513_6273# a_10295_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3897 VPWR ts.ts_ctrl.state\[0\] a_11339_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3898 VGND clknet_0_clk a_8022_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3900 uo_out[0] a_8836_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3901 a_14471_13423# net10 a_14901_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3902 VGND net3 a_16354_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3903 VGND net70 a_16127_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3904 VGND _094_ _111_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3905 VGND a_12313_12234# net21 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3906 a_7929_12015# ts.ts_ctrl.temp_ctr\[8\] a_7847_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3907 VPWR a_16863_1679# a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3908 a_15308_7369# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3910 a_10335_4117# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3911 VPWR a_15123_2197# a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3912 a_17695_4399# a_17507_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3914 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14107_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3915 a_13820_1679# ts.ts_core.dac_vout_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.097 ps=0.975 w=0.65 l=0.15
X3916 VGND a_14347_3615# ts.ts_ctrl.state\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3917 a_11129_9117# _089_ a_11057_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3918 VPWR a_5893_5719# net59 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3919 ts.ts_core.dac_vout_ana_ net14 a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3920 VGND a_3944_14709# _179_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X3921 a_13556_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3922 VGND a_18847_14709# net13 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3924 a_13183_7663# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X3925 a_14935_1941# a_14747_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3926 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3927 VGND _103_ a_12449_9301# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3928 VPWR net60 a_1670_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X3929 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3931 a_14882_7983# _065_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3932 VPWR _109_ a_11150_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3933 VPWR a_16127_5487# a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3934 VGND net69 a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3935 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X3936 VPWR ts.ts_ctrl.temp_ctr\[8\] a_3307_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3937 a_9112_11989# ts.o_res\[7\] a_9934_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3938 VPWR net26 ts.ts_core.capload\[13\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3939 ts.ts_core.dac_vout_ana_ net14 a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3940 VPWR a_17699_13799# a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X3941 a_8459_17759# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3942 VPWR a_7571_1135# a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3943 a_17699_13799# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3944 a_17673_15599# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3945 a_9545_4943# a_9501_5185# a_9379_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3946 VPWR a_11719_2197# a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3947 a_9021_12559# ts.o_res\[15\] a_8583_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3948 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3949 _213_ a_12007_16150# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3950 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3951 a_16315_13103# a_16127_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3952 a_8673_15253# a_8455_15657# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3953 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3954 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3955 VGND ts.ts_ctrl.state\[0\] _112_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3956 a_8590_9295# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
R35 tt_um_hpretl_tt06_tempsens_45.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3957 _147_ a_11467_5825# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X3958 a_6427_16341# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3959 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3960 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3961 a_5140_15253# _190_ a_5269_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3962 a_1769_6895# _160_ a_1551_6807# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3963 VPWR _050_ a_12631_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3964 VPWR _218_ a_8031_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3965 a_15117_11293# _067_ a_15017_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X3966 VGND _093_ a_11931_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3967 a_10689_12559# ts.o_res\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3968 a_7109_18241# a_6891_17999# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3969 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3970 a_15304_7119# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3971 VPWR net70 a_17507_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3972 VPWR a_14571_11623# a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X3973 a_10018_4373# a_9850_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3974 a_8665_12809# _131_ a_8583_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3975 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3976 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3977 a_3763_15823# a_3247_15823# a_3668_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3978 VPWR a_5871_13335# _192_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3979 VGND a_3583_14495# ts.ts_ctrl.temp_ctr\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3980 VPWR a_9524_12559# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3981 a_9353_12809# ts.o_res\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3982 VPWR a_17332_3829# net67 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3983 a_13601_7983# _113_ a_13183_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3984 a_10860_6031# a_9945_6031# a_10513_6273# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3985 net71 a_18243_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3986 a_13183_7663# _122_ _143_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X3987 VPWR a_7263_6879# a_7250_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3988 ts.ts_core.dac_vout_ana_ net71 a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3989 a_14063_10901# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X3990 VPWR a_9245_6005# a_9275_6358# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3991 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3992 VGND _211_ a_9085_18582# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X3993 a_15763_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3994 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3995 VGND a_8619_2223# a_8787_2197# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3996 a_10405_9545# ts.o_res\[5\] a_10321_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3997 a_9128_10159# _087_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3998 a_9188_4943# _007_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3999 VPWR a_10275_4399# a_10443_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4000 a_10275_4399# a_9577_4405# a_10018_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4001 a_16311_4943# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4002 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4003 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4004 a_7565_17999# a_6375_17999# a_7456_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4005 a_5037_10383# a_4993_10625# a_4871_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4006 _098_ a_11606_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4007 VGND net16 a_1633_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4008 a_11991_1941# a_11803_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X4009 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4010 a_12787_7983# _059_ a_12597_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X4011 ts.o_res\[9\] a_12875_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4012 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16499_12821# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4013 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4014 a_14882_7983# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4015 _065_ _059_ a_14471_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4016 a_10138_10927# _088_ a_10138_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X4017 VGND net16 a_4209_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4018 a_13231_12247# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X4019 a_6428_4765# _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4020 a_8300_11247# ts.o_res\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4021 a_18937_2442# ui_in[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4022 a_4135_11231# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4023 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4024 a_16775_7663# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4025 a_6884_6183# ts.ts_ctrl.temp_ctr\[17\] a_7026_6358# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X4026 VPWR a_15483_1135# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4027 a_12332_17833# a_11417_17461# a_11985_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4028 a_10313_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4029 a_7827_17455# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4030 a_11760_14423# ts.o_res\[9\] a_11902_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4031 _054_ _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4032 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4033 VGND net69 a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4034 a_13546_10535# a_13905_10535# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X4035 VPWR clknet_2_1__leaf_clk a_11803_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4037 VPWR a_6651_591# a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4038 a_6741_4373# a_6523_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4039 a_11812_5193# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4040 a_12267_1135# a_12079_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4041 VGND net66 a_6563_16687# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4042 VGND net62 a_3435_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4043 a_4329_13335# a_4425_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X4044 ts.ts_core.capload\[9\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4045 a_10313_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4046 VGND ts.ts_core.dcdel_capnode_ana_ a_5537_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4047 VPWR a_18293_4020# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4048 a_3413_8207# a_3247_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4050 a_10313_2767# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4051 a_11935_16150# a_11753_16150# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4052 VGND net8 a_9792_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X4053 VPWR a_14295_2919# a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X4054 VPWR _212_ a_11343_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R36 net33 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4055 a_10080_9071# _089_ a_9960_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X4056 ts.ts_ctrl.temp_ctr\[4\] a_2111_11231# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X4057 VGND a_13086_11159# _078_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X4058 a_5893_17687# a_5989_17429# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X4059 VGND a_14526_14165# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4060 a_9759_15101# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4061 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12631_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4062 a_16293_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4063 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4064 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4065 VPWR _156_ a_11056_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X4066 uio_out[6] a_12127_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4067 a_1633_12559# a_1589_12801# a_1467_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4068 a_14571_11623# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4069 a_14388_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4070 a_3395_11305# a_2879_10933# a_3300_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4071 VPWR ts.ts_ctrl.state\[1\] a_11435_8864# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R37 tt_um_hpretl_tt06_tempsens_49.LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4072 a_17029_1679# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4073 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_15483_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4074 a_4775_10383# a_4259_10383# a_4680_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4075 a_15308_8457# a_16043_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4076 VPWR a_12547_5095# a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X4077 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4078 _129_ a_7203_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4079 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4080 a_9559_16911# a_9209_16911# a_9464_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4081 VPWR _068_ a_13905_10535# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X4082 VGND net69 a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4083 a_14937_9955# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X4084 a_13733_6941# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.103 ps=1 w=0.42 l=0.15
X4085 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4086 a_16354_9071# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4087 VGND net19 a_7981_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4088 VGND _122_ _143_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4089 VGND a_7815_4917# _211_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4090 a_13845_7369# _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4091 VPWR a_15451_14423# _072_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4092 VGND clknet_2_2__leaf_clk a_2327_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4093 a_14717_9545# _097_ a_14907_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4094 a_11141_3317# a_10975_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4095 VPWR a_9971_743# a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4096 net14 a_17783_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R38 net27 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4097 a_11991_3029# a_11803_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4098 VPWR ts.ts_ctrl.state\[0\] a_10147_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4099 VGND _069_ a_15749_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4100 VGND a_18335_2223# net72 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4101 ts.ts_core.capload\[4\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4102 a_6817_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4103 VPWR _062_ _114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4104 a_10216_14735# a_9135_14735# a_9869_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4105 VGND net70 a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4106 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4107 a_16043_8359# ts.ts_core.dac.vdac_single.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4108 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4109 net67 a_17332_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4110 uo_out[0] a_8836_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4111 a_14471_13423# net10 a_14901_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4112 ts.ts_ctrl.temp_ctr\[13\] a_8459_17759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X4113 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_18755_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4114 _063_ _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4115 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4116 a_12494_17455# a_11417_17461# a_12332_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4117 a_6884_5095# ts.ts_ctrl.temp_ctr\[18\] a_7026_5270# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X4118 a_1585_10383# _165_ a_1367_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4119 ts.ts_core.dac_vout_ana_ net14 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4120 a_11610_8457# _087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4121 a_4972_4777# a_3891_4405# a_4625_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4122 a_7088_4777# a_6007_4405# a_6741_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4123 a_9945_6031# a_9779_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4124 a_9232_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4125 a_16591_1135# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4126 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4127 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4128 a_3247_14735# _172_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X4129 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4130 a_14475_5205# a_14287_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4131 net17 a_6559_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X4132 a_7017_4097# a_6799_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4133 ts.ts_core.dac_vout_ana_ net14 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4134 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4135 VPWR a_16863_2767# a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4136 a_9934_12335# ts.o_res\[7\] a_9112_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4137 uo_out[7] a_9112_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4138 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4139 VGND clknet_2_1__leaf_clk a_9779_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R39 VPWR uio_oe[6] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4140 VGND _205_ a_5363_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4141 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4142 _061_ a_12047_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4143 _133_ a_9597_9955# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X4144 a_14567_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4145 VGND _218_ a_8031_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4146 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4147 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4148 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4149 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12245_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4150 a_17695_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4151 VGND net69 a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4152 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4153 a_6980_13469# _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4154 VPWR a_11975_5461# net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4155 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4156 a_9582_12335# _051_ a_9112_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4157 ts.ts_ctrl.temp_ctr\[6\] a_4411_12319# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4158 a_7539_3829# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4159 VGND net69 a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4160 VGND a_12275_6281# _113_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4161 _014_ _170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4162 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4163 VGND net13 a_15259_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4164 a_11808_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4165 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4166 a_15399_12711# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4167 a_4805_17833# a_3615_17461# a_4696_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4168 a_8877_3829# _153_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X4169 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_16127_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4170 a_7719_15797# ts.ts_ctrl.temp_ctr\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4171 a_8563_15279# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4172 _008_ _159_ a_9865_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4173 VPWR a_10216_14735# a_10391_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4174 a_18937_2442# ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4175 a_16293_13423# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4176 VPWR net13 a_14374_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X4177 a_8679_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4178 a_10331_3671# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X4179 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_15943_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X4180 a_15308_7369# a_16043_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4181 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4182 net1 a_855_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4183 VPWR ts.ts_ctrl.state\[1\] a_16129_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4184 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4185 a_16293_591# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4186 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4187 ts.ts_core.dac_vout_ana_ net14 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4188 VPWR a_15031_4373# a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4189 a_9800_13423# _057_ a_9629_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4190 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4191 a_12320_13897# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X4192 a_15216_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4193 a_14453_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4194 a_18109_10548# _152_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4195 _118_ a_10239_13897# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4196 a_8496_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4197 VPWR a_7815_4917# _211_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4199 ts.o_res\[2\] a_7079_7967# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4200 _029_ a_5455_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4201 VPWR a_4871_17759# ts.ts_ctrl.temp_ctr\[11\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4202 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4203 VPWR a_2111_7093# ts.ts_ctrl.temp_ctr\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4204 VPWR _067_ a_15959_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4205 a_9702_18365# a_9615_18141# a_9298_18251# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X4206 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4207 VGND net67 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4208 VPWR a_8448_15975# _218_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X4209 a_16661_11247# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4210 a_9770_8751# _090_ a_9770_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X4211 ts.ts_ctrl.temp_ctr\[7\] a_4135_11231# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4212 VGND net67 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4214 ts.ts_core.dac_vout_ana_ net14 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4215 a_15465_13647# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4216 a_15216_3017# a_15951_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4217 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4218 VGND net70 a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4219 VPWR net12 a_13546_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X4220 a_12493_7119# _110_ a_12493_7369# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4221 ts.ts_core.dac_vout_ana_ net15 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4222 a_17603_9839# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4223 _048_ a_8532_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X4224 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4225 VPWR a_13967_12711# _088_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4226 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4227 a_14991_14557# net11 a_14900_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X4228 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4229 a_1936_11305# a_855_10933# a_1589_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4231 a_10335_1941# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4232 a_11991_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4233 VPWR _083_ a_7929_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4234 a_11877_15285# a_11711_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4235 VPWR net70 a_16863_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4236 a_8468_10357# _054_ a_9290_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4237 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4238 a_15308_8457# a_16043_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X4239 net18 a_4135_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4240 a_7364_3855# a_6449_3855# a_7017_4097# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4241 a_14707_10901# a_15159_11248# a_15117_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4242 VGND a_9195_15583# a_9129_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4243 VPWR a_8744_5865# a_8919_5791# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4244 a_10493_10159# ts.o_res\[3\] a_10147_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4245 ts.ts_core.dac_vout_ana_ net71 a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4246 a_8774_16406# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X4247 a_7456_17999# a_6541_17999# a_7109_18241# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4248 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16591_10645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4249 a_10299_16885# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4250 a_7827_17455# a_7203_17461# a_7719_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4251 a_13845_7369# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4252 VGND _177_ a_5167_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X4253 a_11124_13897# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X4254 a_12596_5461# a_12447_5540# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4255 a_9283_4943# a_8767_4943# a_9188_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4256 VGND a_4111_4221# a_4279_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4257 VGND a_18293_4020# net5 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4258 ts.ts_core.dac_vout_ana_ net71 a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4259 a_17695_8751# a_17507_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4260 a_10448_11247# _072_ a_10328_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X4261 VGND _212_ a_11343_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4262 a_11991_3029# a_11803_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X4263 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4264 a_8859_13103# _082_ a_9037_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4265 VPWR ui_in[6] a_8399_18543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4266 a_1371_7119# a_1021_7119# a_1276_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4267 a_14545_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4268 a_13901_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4269 VPWR a_4495_16885# _018_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X4270 VPWR a_3299_9269# _164_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4271 _131_ a_7847_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4273 VGND net69 a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4274 VPWR a_2375_12247# _167_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4275 a_13845_7369# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4276 _140_ a_13643_8207# a_14024_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4277 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4278 VPWR a_14379_6575# a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4279 a_12581_4765# a_12537_4373# a_12415_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4280 a_15952_9545# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4281 a_16863_4719# _140_ a_17017_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4282 a_4167_14735# ts.ts_ctrl.temp_ctr\[9\] a_4073_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X4283 a_16293_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4284 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4285 VGND net70 a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4286 ts.ts_core.dac_vout_ana_ net72 a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4287 a_17673_15599# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4288 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4289 a_3013_5853# a_2969_5461# a_2847_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4290 a_4617_6281# ts.ts_ctrl.temp_ctr\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4291 VGND net68 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4292 VPWR a_6559_5487# net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4293 VPWR a_12679_10071# _087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X4294 a_10984_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4295 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4296 a_11056_5193# _155_ a_10965_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X4297 a_3479_6807# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4298 VPWR _065_ _099_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4299 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4300 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4301 VGND a_5423_4917# net16 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4302 net13 a_18847_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4303 VGND a_8399_14735# net19 VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4304 VGND _071_ a_10953_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4305 a_12323_15657# a_11877_15285# a_12227_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4306 VGND a_18937_11636# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4307 VGND _204_ a_5455_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4308 VGND a_17783_5487# net14 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4309 a_11913_16885# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4310 VGND a_4135_11445# net18 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4311 a_9393_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4312 a_6209_8181# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4313 ts.ts_core.dac_vout_ana_ net72 a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4314 ts.ts_core.dac_vout_ana_ net15 a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4315 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4316 a_3413_8207# a_3247_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4317 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4319 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4320 VPWR a_16127_13103# a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X4321 a_8084_5853# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4322 VGND a_7263_9269# a_7197_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4323 a_11521_12809# _117_ a_11425_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4324 a_4956_5461# net59 a_5179_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X4325 a_15487_13909# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4326 VGND a_12875_14709# a_12809_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4327 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4328 a_18671_14451# ui_in[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4329 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4330 a_8632_16599# ts.ts_ctrl.temp_ctr\[11\] a_8774_16406# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X4331 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4332 a_16793_8751# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X4333 VPWR a_11207_7637# uio_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4334 a_5729_14977# a_5511_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4335 a_7088_6953# a_6173_6581# a_6741_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4336 VPWR clknet_2_1__leaf_clk a_8767_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4337 a_12224_4765# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4339 VGND a_10441_5785# a_10375_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4340 VPWR a_10147_3855# a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4341 a_6209_8181# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X4342 VPWR net12 a_14379_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4343 a_15625_14529# net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X4344 a_15308_7369# a_16043_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
R40 VPWR net47 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4345 _065_ _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4346 a_2375_12247# ts.ts_ctrl.temp_ctr\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4347 ts.ts_core.dac_vout_ana_ net14 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4348 VPWR a_9340_11471# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4349 a_7365_15975# a_7461_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X4350 net70 a_17935_13363# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4351 a_2397_15511# a_2493_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X4352 a_6516_11159# ts.ts_ctrl.temp_ctr\[7\] a_6658_10966# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X4353 a_6339_8041# a_5989_7669# a_6244_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4354 a_1573_3855# a_1407_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4355 VPWR a_11913_16885# a_11943_17238# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4356 a_16315_853# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4359 a_14085_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4360 VPWR a_14287_6031# a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4361 VGND _039_ a_10334_18365# VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X4362 VPWR ts.ts_ctrl.state\[0\] a_15591_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4363 VPWR ts.ts_ctrl.state\[0\] a_9687_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X4364 VGND a_12591_11159# _079_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4365 VPWR a_8399_14735# net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4366 a_9524_12559# net8 a_9353_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X4367 a_12892_5603# ts.ts_ctrl.state\[1\] a_12808_5603# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4368 a_4986_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4369 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4370 ts.ts_core.dac_vout_ana_ net14 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4371 a_12591_6895# _112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4372 VPWR clknet_2_1__leaf_clk a_10975_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4373 VGND a_18234_10927# net69 VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X4374 VPWR clknet_2_1__leaf_clk a_13091_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4375 _012_ _167_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4376 VPWR a_16587_7663# a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4378 a_7996_8207# ts.o_res\[18\] a_7775_8534# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X4379 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4380 VGND a_8919_5791# a_8853_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4381 VPWR a_12967_15583# a_12954_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4383 a_3947_4943# a_3431_4943# a_3852_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4384 VPWR a_6833_15253# a_6723_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4385 VPWR a_15535_10357# _094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4386 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4387 _172_ a_3431_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4388 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4389 VPWR a_2014_3967# a_1941_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4390 a_16109_6031# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4392 a_8996_3311# a_8782_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X4393 a_13560_841# a_14295_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4395 a_6427_13621# ts.ts_ctrl.temp_ctr\[11\] a_6825_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X4396 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4397 ts.ts_ctrl.state\[0\] a_12231_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4398 ts.ts_core.dac_vout_ana_ net15 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4399 a_12603_12247# _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4400 ts.ts_ctrl.state\[2\] a_14347_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4401 _086_ a_8859_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X4402 a_14107_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4403 a_13967_12711# a_14331_12533# a_14289_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4404 a_9687_8751# _090_ a_9770_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X4405 a_8496_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4406 a_16960_13647# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4407 a_8782_3311# a_8656_3427# a_8378_3443# VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X4408 VGND _146_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4409 VGND _068_ _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X4410 a_12797_2543# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4411 a_10391_6031# a_9945_6031# a_10295_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4413 a_6251_14709# a_6076_14735# a_6430_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4414 VPWR a_14747_1679# a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X4415 a_12181_7663# _096_ a_11207_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4416 VPWR _143_ a_18325_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4417 VGND a_17935_13363# net70 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4419 a_10335_1941# a_10147_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4421 a_11808_3855# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4422 a_4503_15797# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4423 a_4696_17833# a_3781_17461# a_4349_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4424 a_9091_16406# ts.o_res\[11\] a_8632_16599# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X4425 a_10292_15823# _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4426 VPWR a_16403_1135# a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4427 a_14107_4117# a_13919_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X4428 a_13832_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4429 a_6601_9117# a_6557_8725# a_6435_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4430 _083_ a_14526_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
R41 net31 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4431 a_13755_10429# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X4432 a_16661_11247# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4433 a_5043_11636# _206_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4434 a_17121_7119# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4435 a_6447_7663# a_5823_7669# a_6339_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4436 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4437 a_3570_14191# a_2493_14197# a_3408_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4438 a_10321_13647# ts.ts_ctrl.temp_ctr\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4439 VPWR _071_ a_10229_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4440 a_1573_3855# a_1407_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4441 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_14747_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4442 a_8022_6575# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4443 a_6515_6196# _220_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4444 a_16354_9071# net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4445 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4446 VGND _069_ a_10080_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X4447 VPWR net69 a_16495_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4448 _117_ a_10607_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4449 a_13183_7663# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4450 a_12777_6005# _140_ a_12997_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4451 a_14545_6895# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4452 a_9848_4943# a_8767_4943# a_9501_5185# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4453 a_5423_4917# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4454 VPWR a_16127_5487# a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4455 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4456 a_12819_2223# a_12631_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4457 a_12157_13799# ts.o_res\[13\] a_12320_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4458 VPWR a_7571_1135# a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4459 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4460 a_11851_12247# _066_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X4461 a_15749_10159# _066_ _097_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4462 a_12321_12705# _102_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X4463 ts.ts_ctrl.temp_ctr\[5\] a_2111_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4464 a_11520_7119# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4465 VPWR a_17415_9839# a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4466 VGND net6 a_14882_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4467 VGND a_2111_14709# ts.ts_ctrl.temp_ctr\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4468 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4470 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4472 a_1769_7663# _159_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X4473 a_14901_13423# net10 a_14471_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4474 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4475 ts.ts_core.dac_vout_ana_ net14 a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4476 a_12189_14489# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X4477 _144_ a_12777_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4478 VPWR ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_17507_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4479 a_14907_9545# _097_ a_14717_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X4480 a_11101_11721# _053_ a_11272_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R42 VPWR ts.ts_core.capload\[11\].cap_24.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4481 ts.ts_core.dac_vout_ana_ net72 a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4482 a_15304_7119# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4484 a_1276_14735# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4485 VPWR a_17415_9839# a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4486 a_8877_3829# _153_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4487 a_13992_6031# _063_ a_13769_6296# VGND sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X4488 a_10471_15318# ts.o_res\[14\] a_10012_15511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X4489 a_7847_7663# _090_ a_7929_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4490 VPWR a_8877_9269# a_8907_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4491 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4492 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4493 VPWR _070_ a_12493_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4494 ts.ts_core.dac_vout_ana_ net14 a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4497 a_8455_15657# a_8105_15285# a_8360_15645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4498 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4499 VGND a_9112_11989# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4500 VPWR a_7631_17973# a_7618_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4501 net71 a_18243_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4502 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4503 VGND _107_ a_12449_9301# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4504 a_13327_9813# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X4505 a_9033_591# net33 ts.ts_core.capload\[5\].cap.Y VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4506 VGND _064_ a_14418_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4507 VPWR a_16640_14165# _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4508 VPWR a_9287_3829# _154_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4509 ts.ts_core.dac_vout_ana_ net71 a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4510 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4512 a_10961_13799# ts.o_res\[14\] a_11124_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4513 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4514 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4515 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4516 a_11877_9545# ts.ts_ctrl.temp_ctr\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4517 a_15763_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4518 clknet_2_2__leaf_clk a_4513_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4519 a_18756_15797# uio_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4520 VPWR a_9971_743# a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X4521 a_4621_4943# a_3431_4943# a_4512_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4522 a_2859_5487# a_2235_5493# a_2751_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4523 ts.ts_core.dac_vout_ana_ net15 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4524 a_8958_6358# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X4525 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4526 _059_ net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4527 a_9112_11989# _051_ a_9582_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4528 VGND _171_ a_3431_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X4529 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4530 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref a_16955_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4531 a_8378_3443# a_8656_3427# a_8612_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X4532 a_11991_1941# a_11803_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4533 _059_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X4534 a_13923_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4535 VGND _172_ _014_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4536 VPWR net25 ts.ts_core.capload\[12\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4537 VGND a_5179_16367# _138_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4538 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4539 a_13607_3689# a_13257_3317# a_13512_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4540 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4541 ts.ts_core.dac_vout_ana_ net72 a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4542 VPWR ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_18691_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4543 VGND net70 a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4544 a_6725_13109# a_6559_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4545 a_5619_15101# a_4995_14735# a_5511_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4546 a_9415_1135# a_9227_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4547 a_11877_9545# ts.ts_ctrl.temp_ctr\[1\] a_11793_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4548 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4549 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4550 a_14913_1679# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4551 a_17029_1679# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4552 a_6839_853# a_6651_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4553 a_14085_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4554 a_9245_6005# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X4555 a_4437_8207# a_3247_8207# a_4328_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4556 VPWR a_13643_8207# _140_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R43 net23 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4557 a_4362_5603# _199_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4558 a_18719_5193# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4559 VPWR a_14707_10901# _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X4560 a_6877_15645# a_6833_15253# a_6711_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4561 VPWR _145_ a_15483_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4562 a_4867_12559# a_4517_12559# a_4772_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4563 VPWR net21 a_11325_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4564 a_10952_15823# a_9871_15823# a_10605_16065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4565 VGND _061_ a_14882_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4566 VPWR net11 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4567 ts.ts_ctrl.temp_ctr\[11\] a_4871_17759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4568 a_5094_10966# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X4569 VPWR net12 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4570 a_14085_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4571 a_13183_7663# _122_ _143_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4572 VPWR a_4349_17429# a_4239_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4573 VGND a_12231_3615# a_12165_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4574 a_11417_17461# a_11251_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4575 VPWR net8 a_8415_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4576 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4577 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4578 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9393_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4579 VPWR a_7088_9295# a_7263_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4580 a_16661_11247# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4581 _097_ _066_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4582 VPWR a_6247_5461# a_5989_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X4583 a_16964_13897# a_17699_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4584 a_4073_14735# _172_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4585 VPWR _188_ a_6427_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4586 a_10313_2767# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4587 net18 a_4135_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X4588 a_11724_11247# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4589 a_11593_12809# _116_ a_11521_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4590 _178_ _177_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4591 a_11719_2197# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4592 a_8449_8790# ts.o_res\[3\] a_8235_8790# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X4593 net69 a_18234_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4594 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4595 a_6623_13647# ts.ts_ctrl.temp_ctr\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X4596 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4597 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4598 a_14584_8751# _100_ a_14418_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4599 a_18937_9323# _139_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X4600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4601 a_7981_17821# a_7937_17429# a_7815_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4602 a_17143_14191# a_16955_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4603 a_17695_4399# a_17507_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X4604 a_16591_10645# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4605 a_9020_15657# a_7939_15285# a_8673_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4606 a_11214_6031# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4607 a_13556_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4608 a_17029_1679# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4609 ts.ts_core.dac_vout_ana_ net14 a_16131_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4610 VPWR clknet_2_2__leaf_clk a_4351_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4611 VPWR a_12547_4007# a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4612 a_3859_8207# a_3413_8207# a_3763_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4613 VPWR net2 a_17034_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4614 a_10523_3427# a_10331_3671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X4615 a_9236_841# a_9971_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4616 a_9597_9955# _130_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4617 a_12047_6835# _060_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X4618 a_14500_8751# _097_ a_14584_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4619 _158_ ts.ts_ctrl.temp_ctr\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4620 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13560_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4621 VGND _122_ _143_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4622 VGND _051_ _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4623 a_10359_4399# a_9577_4405# a_10275_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4624 a_11599_3311# a_10975_3317# a_11491_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4625 a_13715_3311# a_13091_3317# a_13607_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4626 a_17121_14511# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4627 net8 a_8399_18543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4629 a_14660_12559# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4630 VGND _085_ a_8859_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4631 net14 a_17783_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4632 VGND a_18335_2223# net72 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4633 VGND a_9800_13423# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4634 a_9800_13423# ts.o_res\[6\] a_9716_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4635 VGND a_8399_14735# net19 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4636 ts.o_res\[17\] a_7263_6879# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4637 VGND a_13546_13335# _082_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X4638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4639 a_4952_11159# ts.ts_ctrl.temp_ctr\[4\] a_5094_10966# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X4640 VGND a_2305_10535# net60 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4641 a_9916_18365# a_9702_18365# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X4642 VPWR a_16127_591# a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4643 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4644 VPWR a_13735_1135# a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X4645 a_7929_7663# ts.ts_ctrl.temp_ctr\[19\] a_7847_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4646 a_12189_14489# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4647 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4648 a_15308_8457# net47 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4649 _154_ a_9287_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X4650 a_10335_3029# a_10147_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4651 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4652 a_1467_11305# a_1021_10933# a_1371_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4653 a_5432_12559# a_4351_12559# a_5085_12801# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4654 _163_ a_2451_9323# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X4655 a_8491_7663# _090_ a_8573_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4656 a_14717_9545# _135_ a_14445_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4657 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4658 ts.ts_core.dac_vout_ana_ net14 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4659 a_6884_6183# ts.o_res\[17\] a_7026_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4660 VPWR _072_ a_12946_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X4661 VPWR a_18937_2442# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4662 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4663 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4664 VPWR _067_ a_13546_10535# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X4665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4666 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4667 VPWR a_17332_3829# net67 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4668 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4669 a_18763_7271# _148_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X4670 a_9025_13103# ts.o_res\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4671 a_14567_12015# a_14379_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4672 a_11977_13103# ts.ts_ctrl.temp_ctr\[13\] a_11895_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4673 a_1589_7361# a_1371_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4674 VPWR a_9020_15657# a_9195_15583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4675 VPWR _065_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4676 ts.ts_core.dac_vout_ana_ net14 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4677 a_15749_8751# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd _134_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4678 a_6880_16911# ts.ts_ctrl.temp_ctr\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X4679 a_5134_4399# a_4057_4405# a_4972_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4680 a_7250_4399# a_6173_4405# a_7088_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4681 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4682 _194_ a_4126_8983# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X4683 VPWR a_12157_9813# _070_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4684 a_7810_17999# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4685 a_14567_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4686 a_14189_9071# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4687 a_9235_1831# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4688 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4689 _211_ a_7815_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4690 VPWR a_9061_16665# a_9091_16406# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4691 a_2014_3967# a_1846_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4692 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4693 uio_out[7] a_14717_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4695 a_6173_6581# a_6007_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4696 a_14664_12809# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4697 VPWR a_16955_8207# a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4698 ts.o_res\[8\] a_5607_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4699 a_9777_17153# a_9559_16911# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4700 _110_ _062_ a_11797_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4701 VPWR ts.ts_ctrl.temp_ctr\[5\] a_2375_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X4702 a_15304_7119# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4703 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4704 a_11672_17821# _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4705 uo_out[4] a_9340_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4706 VPWR ts.o_res\[4\] a_9169_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4707 a_14882_7983# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X4708 VPWR a_14379_12015# a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4709 a_17051_14997# a_16863_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4710 VGND _164_ a_1671_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X4711 VPWR a_8399_14735# net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4712 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4713 a_4993_10625# a_4775_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4714 a_6428_9295# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4715 a_13836_11721# a_14571_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4716 a_12946_13103# _066_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X4717 a_8448_4007# ts.o_res\[19\] a_8590_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4718 a_4713_8751# _192_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X4719 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4720 a_11812_5193# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4721 a_16293_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4722 VPWR a_18671_14451# net9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4723 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4724 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4725 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4726 a_3479_6807# _114_ a_3713_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4727 a_16775_7663# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4728 a_15216_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4729 VPWR a_11045_1367# net57 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4730 a_7829_5493# a_7663_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4731 a_14453_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4732 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4733 a_9615_18141# clknet_2_3__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4734 a_5905_15599# _177_ _188_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4735 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4736 VPWR net30 ts.ts_core.capload\[2\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4737 a_9556_14735# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4738 VPWR a_4993_10625# a_4883_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4739 VGND a_7631_17973# a_7565_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4740 a_11709_3285# a_11491_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4741 ts.o_res\[13\] a_12507_17759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4742 a_3853_7093# ts.ts_ctrl.temp_ctr\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X4743 VPWR a_11272_11471# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4744 a_6185_14735# a_4995_14735# a_6076_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4745 VPWR ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_16955_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4746 net1 a_855_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4747 VPWR a_3571_16586# _017_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4748 a_15216_3017# a_15951_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4749 a_16293_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4750 _169_ _168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4751 ts.ts_core.dac_vout_ana_ net71 a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4752 a_12493_7119# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4753 a_14388_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4754 VGND a_4588_14709# _177_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4755 a_1479_10927# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4756 a_11343_12809# _116_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4757 VGND a_4680_11445# net20 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4759 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _061_ a_16609_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4760 VPWR clknet_2_2__leaf_clk a_6007_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4761 a_15308_8457# a_16043_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4762 VPWR a_12547_5095# a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4763 a_1936_7119# a_1021_7119# a_1589_7361# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4764 a_16661_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4765 VGND net70 a_17029_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4766 VPWR a_18763_7271# _149_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4767 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4768 VPWR a_6904_11471# a_7079_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4769 a_6105_13469# _191_ a_6033_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4771 VPWR _083_ a_7285_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4772 a_14388_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4773 a_7263_9269# a_7088_9295# a_7442_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4774 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4775 VPWR a_10441_15577# a_10471_15318# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4776 a_12596_5461# ts.ts_ctrl.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X4777 VPWR a_11399_1109# a_11141_1109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X4778 a_18756_15797# uio_in[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4779 VPWR a_15031_4373# a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X4780 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4781 VGND clknet_2_2__leaf_clk a_3155_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4782 a_16180_11989# net12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4783 net14 a_17783_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4784 a_11991_3029# a_11803_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4785 a_5909_2543# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4786 VPWR a_5085_12801# a_4975_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4788 a_10313_2767# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4789 VGND net69 a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4791 a_6523_6953# a_6173_6581# a_6428_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4792 VPWR a_16955_7119# a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4793 ts.ts_core.dac_vout_ana_ net15 a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4794 a_13834_8207# _065_ a_14024_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4795 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4796 a_8679_3029# a_8491_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4797 a_8879_4765# a_8625_4438# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X4798 VGND _066_ a_10080_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X4799 a_15952_9545# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4800 a_16293_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4801 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4802 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4803 VPWR a_18848_13621# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4804 VGND a_13059_4703# a_12993_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4805 ts.ts_core.dac_vout_ana_ net72 a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4806 a_3491_11305# a_3045_10933# a_3395_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4807 VGND net68 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4808 a_15304_8207# ts.ts_core.dac.vdac_single.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4809 VGND clknet_2_0__leaf_clk a_5823_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4810 ts.ts_core.dac_vout_ana_ net72 a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4811 VPWR a_6331_12234# _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4812 a_8241_4737# _139_ a_8155_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4813 a_10984_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4814 a_17599_9295# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4815 VGND net10 a_14991_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X4816 a_11325_13103# ts.o_res\[14\] a_11241_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4817 a_5326_4765# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4818 a_1021_7119# a_855_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4819 a_7470_16911# _177_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X4820 a_12875_14709# a_12700_14735# a_13054_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4821 ts.ts_core.capload\[7\].cap.Y ts.ts_core.dcdel_capnode_ana_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4822 a_11679_6183# _112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X4823 a_4871_10383# a_4425_10383# a_4775_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4825 a_12789_13077# ts.o_res\[9\] a_13042_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X4826 a_11610_8457# _122_ a_11518_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X4827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4828 a_9464_16911# _038_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4829 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4830 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.capload\[11\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4831 VGND a_18937_2442# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4832 VGND _074_ a_14937_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0693 ps=0.75 w=0.42 l=0.15
X4833 a_7088_9295# a_6007_9295# a_6741_9537# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4834 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4835 VPWR clknet_2_2__leaf_clk a_5823_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4836 VPWR _164_ a_1775_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X4837 a_9393_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4838 ts.ts_core.dcdel_capnode_ana_ ts.ts_core.i_precharge_n a_13820_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.236 ps=1.38 w=0.65 l=0.15
X4839 VPWR a_4625_4373# a_4515_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4840 VPWR a_6741_4373# a_6631_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4841 VGND net9 a_8456_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X4842 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4843 VGND net19 a_6877_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4844 a_17695_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4845 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4846 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4847 uo_out[1] a_11456_11247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4848 VPWR ts.ts_ctrl.temp_ctr\[4\] a_1585_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4849 a_14475_5205# a_14287_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X4850 VGND _198_ a_4588_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X4851 a_17695_8751# a_17507_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4853 a_7258_8029# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4854 VGND _112_ a_12591_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4855 VGND _068_ a_13905_10535# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X4856 _124_ a_11435_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.26 ps=1.45 w=0.65 l=0.15
X4857 ts.ts_ctrl.temp_ctr\[9\] a_2111_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4858 VPWR ts.ts_ctrl.temp_ctr\[9\] a_2045_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4859 a_13901_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4860 VPWR a_2755_8983# _162_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4861 VGND net38 a_18787_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.236 ps=1.38 w=0.65 l=0.15
X4862 a_11626_16911# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X4863 a_9765_4399# net57 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4864 a_5361_6281# ts.ts_ctrl.temp_ctr\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4865 VPWR a_10147_3855# a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4866 a_17695_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4867 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X4868 a_15948_9295# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4869 a_15308_7369# a_16043_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4870 VPWR clknet_0_clk a_7838_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4871 a_3779_12015# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4872 a_7079_11445# a_6904_11471# a_7258_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4873 _066_ net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4874 a_5780_8359# ts.o_res\[3\] a_5922_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4875 a_15649_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4876 VGND clknet_2_2__leaf_clk a_4351_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4877 VPWR _073_ a_12952_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4878 a_12040_14735# _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4879 ts.ts_core.dac_vout_ana_ net14 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4880 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4881 a_17581_10159# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4882 VGND a_8459_17759# a_8393_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4883 VGND _161_ _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4884 a_8496_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4885 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4886 a_7618_18365# a_6541_17999# a_7456_17999# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4887 a_16315_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4888 VPWR a_14287_6031# a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4889 a_6631_6575# a_6007_6581# a_6523_6953# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4890 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4891 _112_ ts.ts_ctrl.state\[1\] a_15591_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4892 VGND net67 a_11803_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4893 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4894 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4895 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4896 ts.ts_core.dac_vout_ana_ net14 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4897 VPWR a_16587_7663# a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4898 ts.ts_core.dac_vout_ana_ net47 a_15304_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4899 _070_ a_12157_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.38 ps=2.76 w=1 l=0.15
X4900 VGND net67 a_8491_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4901 a_1769_6895# net61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4902 a_10313_3855# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4903 VPWR a_14295_743# a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X4904 VGND _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4905 VGND net67 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4906 _063_ ts.ts_ctrl.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X4907 a_16609_6575# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X4908 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4909 a_5363_15599# _189_ a_5269_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X4910 VPWR a_7355_15583# a_7342_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4912 VGND _080_ a_10977_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X4913 a_3871_8573# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4914 a_9934_12335# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4915 _175_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4918 a_8836_10901# _048_ a_9306_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4919 a_11207_7637# a_11573_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X4920 a_14295_2919# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4921 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4922 ts.ts_core.dac_vout_ana_ net15 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4923 a_11991_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4924 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4925 a_4713_16911# _181_ a_4495_16885# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4927 a_11812_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4928 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4929 _128_ a_10975_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X4930 VPWR net8 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4931 a_6741_6549# a_6523_6953# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4932 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4933 VGND net67 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
R44 VPWR ts.ts_core.capload\[3\].cap_31.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4934 _100_ _099_ a_16127_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X4935 a_14453_6031# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4936 VPWR a_14379_12015# a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4937 a_8496_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4938 a_17143_5205# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4939 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4940 a_7289_15657# a_6099_15285# a_7180_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4941 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4942 _059_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4943 VPWR a_7109_18241# a_6999_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4944 a_12797_2543# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4945 a_12547_743# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4946 a_15535_10357# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4947 a_10335_1941# a_10147_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4948 VGND net69 a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4949 ts.ts_core.dac_vout_ana_ net72 a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4950 VGND net67 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4951 VPWR a_15575_3855# a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X4952 a_1670_10633# _164_ a_1367_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X4953 a_11808_3855# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4954 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4955 VPWR a_17699_13799# a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4956 a_15952_9545# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4957 a_3981_16065# a_3763_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4958 a_14453_6031# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4961 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4962 a_12547_5095# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4963 uo_out[5] a_9524_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4964 VPWR _047_ a_9353_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X4965 VGND net68 a_17029_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
R45 VPWR ts.ts_core.capload\[1\].cap_29.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4966 VPWR a_13546_10535# _090_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X4967 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4968 a_14107_4117# a_13919_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X4969 VPWR clknet_2_3__leaf_clk a_6099_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4970 VPWR a_7815_13407# a_7802_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4971 a_14857_14342# net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X4972 VPWR a_4328_8207# a_4503_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4973 VGND a_10023_4917# a_9957_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4974 a_17121_7119# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4975 VGND a_7079_9055# a_7013_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4976 a_17051_14997# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4977 a_14177_9839# ts.ts_core.i_precharge_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X4978 a_11808_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X4979 a_13183_7663# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4980 a_13280_13423# _081_ a_12789_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X4981 VPWR net69 a_15483_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4982 VGND net17 a_11753_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4983 VPWR a_6559_5487# net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4984 VPWR ui_in[2] a_18278_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4985 a_14347_3615# a_14172_3689# a_14526_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4986 ts.ts_core.dac_vout_ana_ net14 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4988 a_8393_17833# a_7203_17461# a_8284_17833# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4989 a_11045_1367# a_11141_1109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X4990 _202_ a_8879_4438# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X4991 VGND _062_ a_10883_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4992 a_8665_12809# _082_ a_8749_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4993 a_18735_6059# _139_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4995 a_6076_14735# a_5161_14735# a_5729_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4996 _007_ _157_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4997 a_8745_2601# a_7755_2229# a_8619_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4998 VGND _132_ a_9597_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4999 VPWR a_9524_12559# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5000 a_11478_4373# _110_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.136 ps=1.1 w=0.42 l=0.15
X5001 a_9353_12809# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X5002 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X5003 a_13183_7663# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5004 VPWR a_16127_13103# a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5005 a_6515_6196# _220_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5006 VGND a_6883_14887# _186_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5007 a_15741_3855# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5008 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
R46 net24 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5009 VPWR _144_ a_8155_4737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5010 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5011 ts.ts_core.dac_vout_ana_ net71 a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5012 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5013 VPWR a_16127_5487# a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X5014 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5015 VGND clknet_0_clk a_8022_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5017 _105_ a_11711_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X5018 a_11969_1679# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5019 VGND a_11119_4373# _005_ VGND sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.169 ps=1.82 w=0.65 l=0.15
X5020 VGND ts.ts_core.dcdel_capnode_ana_ a_5905_591# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5021 a_5871_13335# ts.ts_ctrl.temp_ctr\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5022 _080_ a_10686_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X5023 net69 a_18234_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5024 a_12397_14735# a_12353_14977# a_12231_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5025 VPWR _083_ a_11977_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5026 a_3944_14709# ts.ts_ctrl.temp_ctr\[8\] a_4167_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X5027 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_13551_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5028 a_3413_15823# a_3247_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5029 a_6515_10058# _219_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5030 a_4239_17455# a_3615_17461# a_4131_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5031 a_6741_9537# a_6523_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5032 uo_out[6] a_9800_13423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X5033 a_9716_13423# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5034 a_2748_14557# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5035 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5036 a_10010_5309# a_8933_4943# a_9848_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5037 VPWR net68 a_16863_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5038 VPWR a_8695_3553# a_8656_3427# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5039 VPWR a_16863_1679# a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X5040 ts.ts_core.dac_vout_ana_ net14 a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5041 a_6447_7663# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5042 a_7045_14735# _184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X5043 VPWR a_15123_2197# a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X5044 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5045 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5046 a_2014_3967# a_1846_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5047 _200_ ts.ts_ctrl.temp_ctr\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5048 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5049 a_16131_6293# a_15943_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5050 VPWR _066_ a_12157_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5051 VPWR a_14379_12015# a_14567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X5052 VPWR _110_ a_12493_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5053 a_10325_14735# a_9135_14735# a_10216_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5054 ts.ts_core.dac_vout_ana_ net14 a_11812_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5055 VPWR _143_ a_18719_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5056 a_5871_13335# ts.ts_ctrl.temp_ctr\[15\] a_6105_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5058 VGND _143_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5059 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5060 _067_ a_16180_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5061 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5062 a_3299_12533# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X5063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5064 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5065 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5066 a_12752_12809# _070_ a_12650_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X5067 a_13821_9117# a_13551_8751# a_13731_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X5068 _113_ a_12275_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X5069 a_14374_13799# a_14843_13621# a_14787_13693# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X5070 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5071 a_9415_1135# a_9227_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X5072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5073 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5074 VPWR a_3853_7093# _195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5075 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5076 _095_ a_14937_9955# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X5077 a_1021_7119# a_855_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5078 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5079 a_11991_1941# a_11803_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5080 VPWR clknet_2_1__leaf_clk net55 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5081 a_13923_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5082 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5083 VPWR a_13555_10901# a_13086_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X5084 a_12862_15101# a_11785_14735# a_12700_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5085 VPWR a_16863_14735# a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5086 VPWR net69 a_16311_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5088 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5089 a_12329_8457# _119_ a_12257_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5090 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5091 _096_ _094_ a_18691_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5092 a_1371_12559# a_1021_12559# a_1276_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5093 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5094 a_7285_12015# ts.ts_ctrl.temp_ctr\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5095 net54 clknet_2_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5096 VPWR a_14571_11623# a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5097 VPWR ts.ts_ctrl.state\[1\] a_11159_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X5098 a_9169_11721# _051_ a_9340_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5099 _091_ a_9770_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X5100 a_14085_3855# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5101 VGND a_9245_6005# a_9179_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5102 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5103 a_11101_11721# ts.o_res\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5104 a_14331_12533# net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5105 a_8782_3311# a_8695_3553# a_8378_3443# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X5106 a_3413_3855# a_3247_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5107 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5108 a_7293_13077# a_7075_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5109 VGND a_11484_17063# _216_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X5110 a_14664_12809# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5111 a_5975_14191# _137_ _190_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X5112 VPWR a_9777_17153# a_9667_17277# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5113 VGND _114_ a_13183_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5114 a_11812_4105# a_12547_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5115 uo_out[2] a_11272_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5116 VPWR net9 a_9277_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X5117 a_13769_6296# _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.209 ps=1.35 w=0.42 l=0.15
X5118 a_12427_4399# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5119 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5120 a_10227_6895# ts.ts_ctrl.temp_ctr\[0\] _158_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5121 a_9460_13799# ts.o_res\[6\] a_9602_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5122 a_3479_6807# _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X5123 a_14882_7983# net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5124 VPWR net7 _140_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5125 a_4425_10383# a_4259_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5126 a_6173_4405# a_6007_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5127 a_4057_4405# a_3891_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5128 _049_ a_8386_11247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X5129 _177_ a_4588_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5130 net72 a_18335_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5131 _095_ a_14937_9955# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.168 ps=1.5 w=1 l=0.15
X5132 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5133 a_13503_10145# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X5134 a_5619_15101# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5135 a_11491_3689# a_10975_3317# a_11396_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5136 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5137 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5138 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5139 a_10495_16189# a_9871_15823# a_10387_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5140 VPWR a_8397_5461# a_8287_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5141 a_2045_7119# a_855_7119# a_1936_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5142 _108_ a_12449_9301# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X5143 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5144 VGND net9 a_9284_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X5145 a_17029_14735# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5146 VGND _064_ a_14471_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5147 a_7079_11445# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5148 a_6934_7446# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X5149 ts.ts_core.dac_vout_ana_ net14 a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5150 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5151 a_17695_4399# a_17507_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5152 _084_ _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5153 VGND a_3413_3311# a_3519_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X5154 VPWR a_16127_5487# a_16315_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5155 a_16354_9071# net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5156 a_11877_15285# a_11711_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5157 a_13556_2767# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5158 a_5537_1455# net31 ts.ts_core.capload\[3\].cap.Y VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5159 VGND net67 a_7571_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5160 a_17673_6895# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5161 a_9393_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5162 VPWR clknet_2_0__leaf_clk net53 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5163 a_11339_6575# a_11159_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5164 a_7155_7119# ts.ts_ctrl.temp_ctr\[2\] a_6792_7271# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5165 _139_ a_12597_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.112 ps=0.995 w=0.65 l=0.15
X5166 a_7640_13481# a_6725_13109# a_7293_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5167 VPWR a_12547_743# a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5168 VPWR _111_ a_13101_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5169 a_6934_7119# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X5170 a_13601_7983# _059_ _143_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5171 a_3576_12381# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5172 a_16569_10383# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5173 a_4513_13621# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5175 _010_ _164_ a_1585_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5176 a_12819_2223# a_12631_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X5177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5178 VGND a_7263_6879# a_7197_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5179 a_13560_841# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5180 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5181 a_4883_10749# a_4259_10383# a_4775_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5182 VGND ts.ts_ctrl.temp_ctr\[12\] _182_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5183 VPWR a_1589_14977# a_1479_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5184 VPWR net9 a_7989_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X5185 net10 a_18848_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5186 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5187 VGND net69 a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5188 VPWR a_17699_13799# a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5189 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd a_18335_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5191 a_11150_9545# _126_ a_11058_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X5192 a_1936_7119# a_855_7119# a_1589_7361# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5193 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5194 a_9941_9295# ts.ts_ctrl.temp_ctr\[0\] a_9503_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5195 VPWR a_8851_3285# a_8782_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X5196 VGND net69 a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5197 VGND a_12231_3615# ts.ts_ctrl.state\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5198 _166_ ts.ts_ctrl.temp_ctr\[4\] a_1858_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X5199 VPWR a_18774_3311# a_18880_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X5200 a_3413_3855# a_3247_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5201 a_11372_11247# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5202 a_15308_8457# net47 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5203 VGND a_7313_4917# a_7247_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5204 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5205 a_6799_3855# a_6449_3855# a_6704_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5206 a_1467_7119# a_1021_7119# a_1371_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5207 VPWR a_15483_11471# a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X5208 a_10335_3029# a_10147_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5209 a_12245_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5210 a_6841_17821# ts.ts_ctrl.temp_ctr\[12\] a_6769_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5211 a_16315_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5212 VGND net9 a_7996_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X5213 a_11793_1455# net36 ts.ts_core.capload\[8\].cap.Y VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5214 VGND _149_ a_13183_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5215 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5216 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5217 VPWR a_9235_1831# a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5218 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5219 a_15649_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5220 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5221 a_4043_4943# a_3597_4943# a_3947_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5222 VGND _073_ a_12952_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X5223 VPWR _027_ a_9414_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X5224 a_7775_8534# ts.o_res\[2\] a_7775_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5225 VGND a_11456_11247# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5226 VGND a_8877_9269# a_8811_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5227 a_10980_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5228 a_16964_13897# a_17699_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X5229 a_4617_6031# _194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
X5230 VPWR a_16187_7895# _060_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X5231 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5233 VPWR a_9287_3829# _154_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5234 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5235 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5236 VGND _067_ a_14011_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5237 a_3491_5791# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5238 a_14567_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5239 a_13836_11721# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5240 a_13595_12336# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5241 a_11895_13103# _082_ a_11977_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5242 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5243 a_8284_17833# a_7369_17461# a_7937_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5244 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5245 VGND _051_ a_11372_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5246 a_15763_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5247 a_13845_7369# _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5248 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15212_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5249 VPWR a_14015_13077# a_13546_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X5250 a_11969_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5251 a_7847_12015# net21 a_7929_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5252 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5253 a_15671_11733# a_15483_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5254 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5255 a_9560_18909# ts.o_res\[12\] a_9339_18582# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5256 a_2401_5493# a_2235_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5257 VPWR _154_ a_8625_4438# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X5258 VPWR a_11719_2197# a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5259 a_16683_10927# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5260 VGND net10 _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5261 a_15304_7119# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5262 ts.ts_ctrl.temp_ctr\[19\] a_5147_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X5263 a_4503_8181# a_4328_8207# a_4682_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5264 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_16127_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5265 a_3395_11305# a_3045_10933# a_3300_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5266 VPWR a_11679_6183# _136_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X5267 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5269 VPWR ts.o_res\[11\] a_9290_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X5270 VPWR net67 a_6651_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5271 VPWR a_15483_1135# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5272 a_12777_6005# net5 a_13079_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X5273 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5274 ts.ts_core.o_tempdelay a_10443_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5275 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5276 VGND _143_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5277 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5278 VPWR a_1936_12559# a_2111_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5279 a_14900_14557# a_14857_14342# a_14828_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X5280 a_4772_12559# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5281 a_16315_13103# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5282 VGND ts.o_res\[13\] a_13280_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5283 VPWR a_18756_15797# net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5284 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5285 uio_out[5] a_14584_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5286 a_11812_5193# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5287 a_12267_1135# a_12079_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5288 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5289 VPWR a_6251_14709# a_6238_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5290 a_13924_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5291 a_17034_9839# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X5292 VGND _061_ a_14882_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5293 a_14453_6031# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5294 a_8481_7369# ts.ts_ctrl.temp_ctr\[18\] a_8399_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5295 VGND net17 a_12581_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5296 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5297 a_14583_13693# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X5298 a_17029_14735# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5299 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5300 a_10313_2767# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5301 a_12691_7663# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X5302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5303 a_16298_4719# net65 a_16129_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X5304 VPWR a_16863_2767# a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X5305 a_4156_7119# ts.ts_ctrl.state\[2\] a_3853_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5306 ts.ts_ctrl.temp_ctr\[0\] a_10023_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X5307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5308 a_2751_15253# ts.ts_ctrl.temp_ctr\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5309 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5310 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5311 a_16127_10159# _095_ _100_ VGND sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X5312 VGND a_6059_6005# _137_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5313 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5314 a_13086_11159# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X5315 VGND net19 a_12397_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5316 a_6907_4221# a_6283_3855# a_6799_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5317 uio_out[6] a_12127_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5318 a_16793_8751# _061_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5319 a_11255_4399# ts.ts_ctrl.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5321 VGND net70 a_14660_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5322 VPWR _083_ a_10321_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5323 a_10216_14735# a_9301_14735# a_9869_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5324 a_2843_14569# a_2327_14197# a_2748_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5325 a_14388_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5326 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5327 a_8109_2223# ts.ts_core.tempdelay_async VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5328 VGND net17 a_8413_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X5329 VPWR ts.ts_ctrl.state\[1\] a_13731_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5330 a_2659_10357# ts.ts_ctrl.temp_ctr\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5331 a_9306_11247# _049_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X5332 a_8614_11721# ts.o_res\[16\] a_8532_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5333 a_14913_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5334 VPWR a_16955_8207# a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5335 a_14857_10383# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X5336 _085_ a_7847_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5337 VGND ts.ts_ctrl.temp_ctr\[15\] _189_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5338 a_7079_9055# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5339 a_10677_9295# ts.o_res\[1\] a_10239_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5340 VPWR ts.ts_ctrl.state\[0\] _156_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5341 _050_ net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5342 a_14707_10901# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.143 ps=1.33 w=0.42 l=0.15
X5343 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_15483_1135# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5344 a_15308_8457# a_16043_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5345 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5346 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5347 a_13560_3017# a_14295_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5348 net56 a_3519_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X5349 a_14567_12015# a_14379_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5350 _059_ net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X5351 a_10605_16065# a_10387_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
R47 VPWR ts.ts_core.capload\[5\].cap_33.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5352 a_14445_9545# _134_ a_14195_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5353 VGND a_3571_16586# _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5354 VGND a_18243_1135# net71 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5355 a_16477_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5356 a_6331_12234# _209_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5357 a_15315_10383# _067_ a_15125_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5358 a_9415_2223# a_9227_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5359 VGND _066_ a_10448_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X5360 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9415_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5361 a_6185_1679# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5362 a_17029_2767# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5363 a_16609_6575# _061_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5364 a_15216_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5365 a_7921_2229# a_7755_2229# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5366 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5367 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5368 a_6817_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5369 a_9919_13974# ts.o_res\[6\] a_9460_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X5370 a_11991_3029# a_11803_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5371 ts.ts_core.i_precharge_n a_13705_6353# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.146 ps=1.34 w=1 l=0.15
X5372 VPWR _062_ _114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5373 a_12231_3615# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5374 VPWR a_16127_13103# a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5375 VGND a_13611_4917# net68 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X5376 a_14664_12809# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5377 a_10313_2767# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5378 VGND net69 a_17673_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5379 a_15487_13909# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5380 VPWR ts.ts_core.dac_vout_ana_ a_13643_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.321 pd=1.68 as=0.109 ps=1.36 w=0.42 l=0.15
X5381 a_8744_5865# a_7829_5493# a_8397_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5382 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5383 ts.ts_core.dac_vout_ana_ net15 a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5384 VGND _047_ a_9658_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5385 ts.ts_core.dac_vout_ana_ net14 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5387 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5388 VPWR a_7079_7967# a_7066_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5389 a_8877_9269# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5390 a_7197_4777# a_6007_4405# a_7088_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5391 VPWR _143_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5392 VGND a_2111_9055# a_2045_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5393 a_13836_11721# a_14571_11623# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X5394 a_17121_14511# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5395 ts.ts_ctrl.temp_ctr\[15\] a_6251_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X5396 VPWR a_6651_591# a_6839_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5397 a_15304_8207# ts.ts_core.dac.vdac_single.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5398 VGND a_9889_13621# a_9823_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5399 a_5085_12801# a_4867_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5400 a_16964_13897# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5401 VGND a_6247_17429# a_5989_17429# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X5402 a_10984_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5403 a_10147_9839# _069_ a_10229_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5404 VPWR net12 a_14733_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X5405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5406 a_10335_1941# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5407 a_8749_12809# ts.ts_ctrl.temp_ctr\[15\] a_8665_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5409 VGND a_8022_6575# clknet_2_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5410 VPWR a_13735_1135# a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5411 VPWR ts.o_res\[5\] a_9353_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5413 a_16315_13103# a_16127_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5414 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5415 a_12319_4777# a_11803_4405# a_12224_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5416 net69 a_18234_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5417 a_14545_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5419 a_14567_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5420 a_9524_12559# _056_ a_9353_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5421 a_9020_15657# a_8105_15285# a_8673_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5422 VPWR a_17332_3829# net67 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5423 VPWR a_16127_2223# a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5424 _141_ a_16465_5193# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.373 ps=1.75 w=1 l=0.15
R48 VPWR ts.ts_core.capload\[4\].cap_32.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5425 a_17695_6575# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5426 ts.ts_core.capload\[9\].cap.Y net37 a_6277_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5427 VGND _106_ a_10239_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5428 VGND clknet_2_0__leaf_clk a_3431_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5429 a_15017_11293# _068_ a_14928_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0619 ps=0.715 w=0.42 l=0.15
X5430 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5431 _074_ a_17191_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5432 VGND clknet_2_2__leaf_clk a_3247_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5433 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5434 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5435 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5436 a_10124_16911# a_9209_16911# a_9777_17153# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5437 a_6704_3855# _046_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5438 a_13901_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5439 a_1589_14977# a_1371_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5440 a_7250_9661# a_6173_9295# a_7088_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5441 a_6741_9537# a_6523_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5442 VPWR a_16955_7119# a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5444 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5445 VPWR a_10147_3855# a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X5446 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5447 a_6449_3855# a_6283_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5448 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5449 a_15948_9295# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5450 a_11711_9295# _087_ a_11889_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5451 a_7534_15645# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5452 a_15308_7369# a_16043_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5453 a_13327_9813# a_13503_10145# a_13455_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X5454 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5455 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5456 a_1276_11293# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5457 VGND _111_ a_12851_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5458 a_6619_4777# a_6173_4405# a_6523_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5459 a_13603_12533# net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X5460 VPWR a_3960_11305# a_4135_11231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5461 ts.ts_core.dac_vout_ana_ net14 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5462 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5463 VPWR a_9869_14977# a_9759_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5464 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X5465 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5466 VPWR _081_ a_9025_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X5467 a_16960_13647# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5468 VGND _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5469 VGND net67 a_8657_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5470 a_7343_6358# ts.o_res\[17\] a_6884_6183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X5471 a_16315_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5472 uio_out[4] a_11207_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5473 net18 a_4135_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5474 VPWR net19 a_9916_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X5475 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5476 _125_ a_12079_8457# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X5477 a_10037_15823# a_9871_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5478 ts.ts_core.dac_vout_ana_ net14 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5479 VGND net17 a_6601_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5480 VPWR _137_ a_5179_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5481 ts.ts_core.dac_vout_ana_ net14 a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5482 _023_ _194_ a_3701_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5483 a_7153_17999# a_7109_18241# a_6987_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5484 a_15216_3017# a_15951_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5485 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5486 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5487 VPWR a_13059_4703# a_13046_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5488 a_2751_5865# a_2235_5493# a_2656_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5489 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5490 VPWR net69 a_17507_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5491 VPWR a_12591_11159# _079_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5492 ts.ts_core.dac_vout_ana_ net14 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5493 a_2957_10205# _159_ a_2869_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X5494 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5495 a_2751_6549# ts.ts_ctrl.temp_ctr\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5496 a_7079_9055# a_6904_9129# a_7258_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5497 VPWR a_2439_4123# a_2355_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5498 VPWR _064_ _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5499 a_17603_9839# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5500 VGND ui_in[6] a_8399_18543# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X5501 VPWR a_3491_5791# a_3478_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5502 a_13556_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5503 a_16298_4719# ts.ts_ctrl.state\[0\] a_16212_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X5504 a_14296_4399# a_15031_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X5505 VGND clknet_2_2__leaf_clk a_855_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5506 _114_ _062_ a_12591_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5507 a_17599_9295# _140_ a_17753_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5508 a_11812_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5509 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5511 _122_ _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5512 VGND a_7286_9839# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5513 a_9232_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5514 a_11812_841# a_12547_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X5515 a_10154_15645# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X5516 a_6833_15253# a_6615_15657# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5517 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9227_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5518 a_16315_853# a_16127_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5519 a_13455_10205# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X5520 VPWR rst_n a_855_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5521 _109_ a_11339_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X5522 VGND a_18763_9447# _152_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5524 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd _065_ a_16771_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5525 a_11053_5719# ts.ts_core.o_tempdelay VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X5526 VGND _174_ _015_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5527 VPWR _099_ a_18763_9447# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5528 a_9957_4943# a_8767_4943# a_9848_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5529 _171_ a_2787_10205# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X5530 a_15671_11733# a_15483_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5531 a_9340_11471# ts.o_res\[12\] a_9169_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X5532 VPWR a_16687_9447# a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5533 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5534 ts.ts_core.dac_vout_ana_ net15 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5535 VPWR _204_ a_5455_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5536 a_17029_2767# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5537 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _061_ a_16609_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5538 VPWR _051_ a_11101_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X5539 VPWR _072_ a_11851_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5540 a_11991_3029# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5541 ts.ts_core.dac_vout_ana_ net72 a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5542 a_6796_17999# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
R49 ts.ts_core.capload\[15\].cap_28.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5543 VGND a_7631_17973# ts.ts_ctrl.temp_ctr\[12\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5544 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.capload\[5\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5545 a_14453_6031# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5546 a_2111_14709# a_1936_14735# a_2290_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5547 _062_ ts.ts_ctrl.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5548 a_1021_12559# a_855_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5549 a_11272_11471# _050_ a_11101_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X5550 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5551 a_3944_14709# ts.ts_ctrl.temp_ctr\[10\] a_4073_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X5552 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14287_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5553 a_16293_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5555 VGND a_6251_14709# a_6185_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5556 a_14717_9545# _138_ a_14195_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5557 VPWR a_6515_5108# _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5558 a_11808_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5559 a_6839_853# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5560 a_11338_4719# _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.258 ps=1.45 w=0.65 l=0.15
X5561 net70 a_17935_13363# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X5562 a_10403_6397# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5563 a_16293_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5564 a_6904_11471# a_5823_11471# a_6557_11713# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5565 VPWR a_4135_11445# net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X5566 a_11337_13423# ts.o_res\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5567 a_6449_3855# a_6283_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5568 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5569 uo_out[7] a_9112_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5570 a_18671_14451# ui_in[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X5571 a_11417_17461# a_11251_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5572 a_16293_591# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5573 ts.ts_ctrl.state\[1\] a_13059_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5574 a_3481_13675# _172_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X5575 VPWR _114_ a_12691_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X5576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5577 VGND net12 a_14379_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5578 a_16293_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5579 _075_ a_14707_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X5580 VPWR a_15465_3311# a_15571_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5582 a_11101_11721# _050_ a_11272_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5583 VPWR a_12507_17759# a_12494_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5584 a_6891_17999# a_6375_17999# a_6796_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5585 VPWR a_11053_5719# _153_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X5586 a_13540_5487# _140_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X5587 VGND ts.ts_ctrl.temp_ctr\[6\] a_2849_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5588 VPWR net19 a_9095_17973# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5589 ts.ts_core.dac_vout_ana_ net72 a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5590 a_9393_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5591 VGND net67 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5592 _123_ a_8399_7369# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5593 ts.ts_core.dac_vout_ana_ net15 a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5594 a_7343_5270# ts.o_res\[18\] a_6884_5095# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X5595 _174_ _114_ a_3247_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5596 a_5905_591# net22 ts.ts_core.capload\[0\].cap.Y VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5597 VGND a_2751_6549# a_2493_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X5598 a_9195_15583# a_9020_15657# a_9374_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5599 VPWR clknet_2_0__leaf_clk a_5823_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5600 VGND net4 a_18597_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5601 VPWR a_8673_15253# a_8563_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5603 net68 a_13611_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X5604 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10147_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5605 VGND _047_ a_9934_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5606 VGND a_9112_11989# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X5607 VPWR ts.ts_ctrl.temp_ctr\[18\] a_4617_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5608 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5609 a_11035_6005# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5610 ts.ts_core.dac_vout_ana_ net14 a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5611 net17 a_6559_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5612 _127_ a_10138_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X5613 VGND clknet_2_3__leaf_clk a_6559_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5614 a_11812_4105# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5615 ts.ts_core.dac_vout_ana_ net71 a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5617 VPWR clknet_2_2__leaf_clk a_855_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5618 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5619 VPWR a_6741_9537# a_6631_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5620 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5621 VPWR a_12231_3615# a_12218_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5622 a_5411_10966# ts.o_res\[4\] a_4952_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X5623 VPWR a_10147_3855# a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5624 VPWR a_12157_13799# _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X5625 a_11216_5603# ts.ts_core.o_tempdelay VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X5626 a_9667_17277# a_9043_16911# a_9559_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5627 VPWR a_1936_7119# a_2111_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5628 a_17695_8751# a_17507_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X5629 a_1021_8757# a_855_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5630 VGND ts.o_res\[15\] a_9582_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5631 a_10759_7119# ts.ts_ctrl.temp_ctr\[0\] a_10668_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X5632 a_3300_11293# _014_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5633 a_14107_4117# a_13919_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5634 a_13832_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5635 VPWR a_7159_16599# _184_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X5636 a_15304_8207# net47 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5637 VPWR _139_ a_18763_8359# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5638 a_13231_12247# a_13595_12336# a_13553_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5639 VGND _138_ _014_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5640 a_5085_12801# a_4867_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5641 VPWR clknet_2_3__leaf_clk a_11251_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5642 ts.ts_core.dac_vout_ana_ net14 a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5643 VPWR a_14379_6575# a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5644 VGND net7 a_11606_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X5645 a_11573_7663# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5646 VPWR net8 a_8614_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5647 VGND net67 a_15943_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5648 VGND a_8459_17759# ts.ts_ctrl.temp_ctr\[13\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5650 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5651 a_16131_6293# a_15943_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5652 a_17603_9839# a_17415_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5653 a_3781_17461# a_3615_17461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5654 VPWR a_12127_7093# uio_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5655 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5656 a_15649_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5657 VGND _143_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5658 VPWR net13 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5659 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5660 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5661 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X5662 VPWR a_13595_12336# a_13231_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X5663 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5664 a_13463_5807# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5665 a_11484_17063# ts.o_res\[13\] a_11626_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5666 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5667 a_11696_8207# ts.ts_ctrl.temp_ctr\[2\] a_11435_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5668 VPWR a_8468_10357# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5669 _040_ a_10975_17455# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5670 a_11969_1679# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5671 a_10321_13897# ts.ts_ctrl.temp_ctr\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5672 a_8194_2223# a_7755_2229# a_8109_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5673 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5674 a_11724_11247# _052_ a_11456_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5675 VPWR a_16495_10927# a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5676 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5677 a_7365_15975# a_7461_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X5678 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5679 a_10932_10633# _076_ a_10830_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X5680 a_9290_10633# _054_ a_8468_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5682 a_12789_13077# _081_ a_12946_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X5683 VGND net67 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5684 VPWR net27 ts.ts_core.capload\[14\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5685 a_1479_15101# a_855_14735# a_1371_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5686 a_5893_5719# a_5989_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X5687 a_5085_5807# _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X5688 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5689 a_8496_1679# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5690 net11 a_18756_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5691 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5693 ts.ts_core.capload\[11\].cap.Y net24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5694 a_11573_7663# _070_ a_11573_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5695 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5696 a_12797_2543# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5697 a_16591_10645# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5698 a_1276_7119# _009_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5699 VPWR a_5043_11636# _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5700 a_10335_1941# a_10147_1679# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X5701 a_13560_841# a_14295_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X5702 ts.ts_core.dac_vout_ana_ net72 a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5703 VGND net67 a_16403_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5704 a_18848_13621# uio_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5705 a_2045_14191# _173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X5706 a_7263_6879# a_7088_6953# a_7442_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5707 a_3763_15823# a_3413_15823# a_3668_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5708 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5709 a_10557_6031# a_10513_6273# a_10391_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5710 a_8590_15823# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X5711 _041_ a_9595_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5712 a_17143_5205# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5713 VGND net8 a_10068_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X5714 a_11812_4105# a_12547_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5715 VGND _114_ a_13183_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5716 _073_ a_16640_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5717 a_11985_17429# a_11767_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5718 a_9945_4399# a_9411_4405# a_9850_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5719 VPWR ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_17332_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5720 a_6101_17161# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5721 VGND _081_ a_9021_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X5722 a_16960_13647# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5723 a_15465_3311# a_15229_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X5724 a_7829_5493# a_7663_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5725 VPWR _159_ a_1775_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X5726 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5727 VPWR a_15575_3855# a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5728 VGND net68 a_17507_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5729 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15948_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5730 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5731 a_11808_4943# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5732 a_9770_8751# ts.ts_ctrl.temp_ctr\[16\] a_9687_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5733 a_14660_12559# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5734 a_8991_8534# a_8809_8534# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5735 VGND a_9800_13423# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5736 VGND a_18847_16341# net12 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5737 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5738 _189_ ts.ts_ctrl.temp_ctr\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5739 a_15487_13909# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5740 VPWR _184_ _185_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5741 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5742 VGND net67 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5743 a_2397_6807# a_2493_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X5744 a_17121_7119# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5745 VPWR _065_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5747 a_17673_9071# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5748 VPWR net69 a_14379_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5749 _132_ a_8583_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5750 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5751 a_12161_8457# _124_ a_12079_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X5752 a_10375_15645# ts.ts_ctrl.temp_ctr\[14\] a_10012_15511# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5753 a_11812_841# a_12547_743# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5754 VPWR net23 ts.ts_core.capload\[10\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5755 a_9415_1135# a_9227_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5757 a_15125_10383# _067_ a_15315_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5758 VGND a_6515_5108# _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
R50 net22 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5759 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5760 a_12797_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5761 VPWR a_14015_10357# a_13546_10535# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X5762 VGND a_13059_4703# ts.ts_ctrl.state\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5763 a_8811_3855# ts.ts_ctrl.temp_ctr\[19\] a_8448_4007# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5764 VPWR _169_ a_3299_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X5765 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5766 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5767 a_18847_14709# uio_in[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X5768 VPWR a_4972_4777# a_5147_4703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5769 a_8320_2601# a_7921_2229# a_8194_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5771 VPWR a_9340_11471# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5772 a_9169_11721# ts.o_res\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5773 VGND a_7838_14191# clknet_2_3__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5774 VGND ts.ts_ctrl.temp_ctr\[7\] _170_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5775 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5776 a_12127_7093# _125_ a_13101_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5777 VPWR ts.ts_ctrl.temp_ctr\[1\] a_10294_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X5778 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5779 VGND a_2397_15511# net64 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5780 a_9063_8534# ts.o_res\[1\] a_9063_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5781 a_15535_10357# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5782 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5783 VPWR a_14747_1679# a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5784 a_9658_11247# ts.o_res\[0\] a_8836_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5785 a_17121_14511# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5786 a_10495_16189# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5787 a_15451_14423# net12 a_15625_14529# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5788 a_10953_12559# ts.o_res\[2\] a_10607_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5789 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5790 a_8717_15645# a_8673_15253# a_8551_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5791 a_11808_4943# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5792 a_3597_4943# a_3431_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5793 VGND net70 a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X5794 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5795 a_15671_11733# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5796 a_14177_9839# a_14011_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X5797 a_7703_8534# a_7521_8534# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5798 a_12132_15645# _037_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5799 a_17695_15279# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5800 VGND a_12231_3615# ts.ts_ctrl.state\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5801 VPWR ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_17783_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5802 VGND _129_ a_9214_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X5803 VPWR a_13231_12247# _081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5804 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5805 a_1021_12559# a_855_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5806 a_6523_6953# a_6007_6581# a_6428_6941# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5807 a_11061_15823# a_9871_15823# a_10952_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5808 a_4328_15823# a_3247_15823# a_3981_16065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5810 a_12357_6281# _112_ a_12275_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5811 a_12245_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5812 a_10860_6031# a_9779_6031# a_10513_6273# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5813 a_7286_9839# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5814 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref _148_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5815 VPWR a_8175_3285# ts.o_res\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X5816 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref a_17121_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5817 a_12631_8457# _059_ _122_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5818 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X5819 a_9353_12809# _056_ a_9524_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5820 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5821 a_11931_7983# _093_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5822 VGND a_14374_13799# _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X5823 VGND a_14347_3615# ts.ts_ctrl.state\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5824 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5825 VPWR a_11035_6005# a_11022_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5826 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5827 VGND net16 a_1633_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5828 VGND net9 a_8386_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X5829 ts.ts_core.dac_vout_ana_ net15 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5830 VGND a_6559_5487# net17 VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X5831 a_16964_13897# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5833 VGND net9 _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5834 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13928_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5835 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5836 a_6382_12886# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X5837 a_13601_7983# _059_ _143_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5838 a_8275_5865# a_7829_5493# a_8179_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5839 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5840 a_1589_7361# a_1371_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5841 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5842 a_4312_4765# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5843 VPWR a_11719_2197# a_10984_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5844 _154_ a_9287_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5845 a_3316_5865# a_2401_5493# a_2969_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5847 a_1861_13103# _166_ a_1777_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5848 a_13923_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5849 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5850 a_17681_9545# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5851 _107_ a_10239_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5852 net18 a_4135_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5853 a_6382_12559# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X5854 a_13832_11471# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5855 a_6983_15797# ts.ts_ctrl.temp_ctr\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5856 VPWR net68 a_14287_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5857 VGND a_10391_14709# a_10325_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5858 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15741_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5859 VPWR a_9501_5185# a_9391_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5860 VGND net16 a_4025_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5861 uio_out[5] a_14584_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5862 VGND ts.ts_ctrl.temp_ctr\[3\] _161_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5863 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_11969_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5864 a_11517_4943# _062_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5866 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5867 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5868 VPWR a_4328_15823# a_4503_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5869 a_11241_13103# _120_ a_11159_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5870 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5871 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5872 _138_ a_5179_16367# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5873 a_2045_14735# a_855_14735# a_1936_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5874 a_16361_8001# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X5875 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5876 VPWR a_11851_12247# _116_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X5877 VPWR a_3307_13799# _173_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X5878 res1_n a_2439_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5879 a_2111_7093# a_1936_7119# a_2290_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5880 VPWR a_5381_11225# a_5411_10966# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5881 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5882 a_18243_7983# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5883 a_14584_8751# _108_ a_14418_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5884 a_12673_12015# a_12603_12247# _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
X5885 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5886 VPWR a_3583_14495# a_3570_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5887 a_4075_6031# ts.ts_ctrl.temp_ctr\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5888 _015_ _173_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5889 VPWR a_8491_2767# a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5890 VPWR a_15483_11471# a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5892 VPWR a_16955_8207# a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5893 a_8703_2223# a_7921_2229# a_8619_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5894 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
R51 uio_oe[1] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5895 VGND _194_ a_4156_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5896 VPWR _211_ a_9085_18582# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X5897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5898 a_17029_2767# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5899 VGND a_6884_6183# _220_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X5900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5901 _041_ a_9595_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5902 a_6240_12711# ts.ts_ctrl.temp_ctr\[8\] a_6382_12886# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5903 ts.ts_ctrl.temp_ctr\[12\] a_7631_17973# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X5904 a_13560_3017# a_14295_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5906 net8 a_8399_18543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X5907 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.capload\[15\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5908 ts.ts_core.dac_vout_ana_ net15 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5909 _065_ _059_ a_14471_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5910 _055_ a_8235_8790# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X5911 VGND _078_ a_12809_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X5912 a_4669_4765# a_4625_4373# a_4503_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5913 VPWR _133_ a_14195_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5914 a_6785_4765# a_6741_4373# a_6619_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5915 VGND a_18243_1135# net71 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5917 _104_ a_11435_8864# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X5918 a_7197_9295# a_6007_9295# a_7088_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5919 a_9577_4405# a_9411_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5921 a_13054_14735# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5922 a_5179_5807# _200_ a_5085_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5923 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5924 VPWR a_12792_15657# a_12967_15583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5925 a_9759_15101# a_9135_14735# a_9651_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5926 a_14384_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X5927 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5928 a_17029_2767# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5929 a_10375_5853# _058_ a_10012_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5930 a_15216_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5931 VPWR a_13603_12533# _068_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5932 a_1467_12559# a_1021_12559# a_1371_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5933 a_3981_16065# a_3763_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5934 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_15943_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5935 VGND net20 a_10649_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5936 VPWR _065_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5937 VGND a_17332_3829# net67 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5938 ts.ts_ctrl.temp_ctr\[9\] a_2111_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5939 a_5989_7669# a_5823_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5940 a_8811_15823# ts.ts_ctrl.temp_ctr\[15\] a_8448_15975# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X5941 VGND a_7539_3829# a_7473_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5942 a_14289_12559# net13 a_14189_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X5943 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_13901_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X5944 a_17034_9839# _061_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5945 _144_ a_12777_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5946 a_15308_8457# net47 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5947 a_11272_11471# _053_ a_11101_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5948 VGND a_8448_15975# _218_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X5949 a_10335_3029# a_10147_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X5950 VPWR _143_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5951 VGND clknet_2_3__leaf_clk a_6099_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5952 a_14664_12809# a_15399_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5953 a_10335_1941# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5954 VPWR a_17783_5487# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5955 a_12851_7119# a_12493_7369# a_12127_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5956 a_7342_15279# a_6265_15285# a_7180_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5957 a_7258_11471# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5958 a_6428_4765# _045_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5959 a_10977_9955# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5960 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5961 a_9913_14735# a_9869_14977# a_9747_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5962 ts.ts_core.dac_vout_ana_ net71 a_10335_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X5963 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5964 a_1371_9129# a_855_8757# a_1276_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5965 VGND net18 a_5129_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5968 a_4259_14557# ts.ts_ctrl.temp_ctr\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5969 VPWR a_16127_2223# a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5970 a_6619_9295# a_6173_9295# a_6523_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5971 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5972 a_6980_13469# _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
R52 tt_um_hpretl_tt06_tempsens_41.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5973 clknet_2_1__leaf_clk a_8022_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5974 a_10328_11247# ts.o_res\[11\] a_10138_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X5975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5976 VPWR net11 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5977 a_17673_15599# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5978 a_15304_7119# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5979 VPWR clknet_2_0__leaf_clk a_855_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5980 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5981 a_9643_14410# _208_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5982 VPWR a_16955_7119# a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X5983 a_6883_14887# _184_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X5984 a_13832_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5985 a_3852_4943# _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5986 a_16661_11247# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5987 a_4495_16885# _181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X5988 VPWR net70 a_16955_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5989 VGND _104_ a_11711_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5990 _160_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5991 ts.ts_core.dac_vout_ana_ net72 a_14384_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5992 VPWR _171_ a_3431_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5993 _176_ a_4259_14557# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X5994 VGND net18 a_1633_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5995 a_12245_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5996 a_10295_6031# a_9779_6031# a_10200_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5997 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5998 a_15304_8207# ts.ts_core.dac.vdac_single.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5999 VGND net4 a_16170_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6000 a_7838_14191# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6001 a_10984_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6002 VGND a_8448_9447# _219_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X6003 a_10596_7119# a_10147_7119# a_10294_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6004 VPWR clknet_2_2__leaf_clk a_3615_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6005 a_9112_11989# ts.o_res\[15\] a_9500_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6006 VPWR a_13735_1135# a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6007 _059_ net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6008 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6009 a_12245_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6010 ts.ts_core.dac_vout_ana_ net14 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6011 VPWR a_12547_743# a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6012 VGND clknet_2_2__leaf_clk a_2879_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X6014 a_8415_13103# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6015 a_8590_16150# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X6016 a_1677_14511# _175_ a_1459_14423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6017 ts.ts_core.dac_vout_ana_ net14 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6018 VPWR a_16127_591# a_16315_853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6019 a_3617_8751# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6020 uo_out[3] a_8468_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6021 a_8563_15279# a_7939_15285# a_8455_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6022 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6023 ts.ts_core.dac_vout_ana_ net15 a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6024 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6025 ts.ts_core.dac_vout_ana_ net71 a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6026 a_1936_12559# a_855_12559# a_1589_12801# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6027 a_9415_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6028 a_14195_9295# _138_ a_14717_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6029 VPWR _100_ a_14852_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6030 _120_ a_10975_8864# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6031 a_11456_11247# _052_ a_11724_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6032 _114_ _062_ a_12591_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6033 a_13555_10901# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X6034 VGND _177_ _178_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6035 _122_ _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6036 VPWR a_14843_13621# a_14374_13799# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6037 a_16775_7663# a_16587_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6038 VPWR a_12587_15988# _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6039 a_2755_8983# ts.ts_ctrl.temp_ctr\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6040 a_8938_10633# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6041 VPWR net13 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6042 VGND net19 a_8717_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6043 a_9751_9955# _130_ a_9679_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6044 VGND a_12789_13077# _101_ VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X6045 a_9821_16911# a_9777_17153# a_9655_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6046 a_12587_15988# _213_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6047 ts.o_res\[18\] a_7263_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6048 VPWR a_16687_9447# a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X6049 _096_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd a_18243_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6050 VPWR _067_ a_14063_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X6051 net52 clknet_2_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6052 a_17141_4399# net2 a_17017_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.235 ps=1.47 w=1 l=0.15
X6053 a_13825_3285# a_13607_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6054 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6055 a_6792_7271# ts.o_res\[2\] a_6934_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6056 a_19057_3311# a_18880_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X6057 ts.ts_core.dac_vout_ana_ net72 a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6058 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6059 a_10686_10383# _079_ a_10932_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X6060 VGND _128_ a_9597_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6061 VPWR a_18109_10548# ts.ts_core.dac.vdac_single.en_pupd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6062 a_14453_6031# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6064 a_10313_2767# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6065 VGND rst_n a_855_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6066 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6067 a_6603_12559# ts.ts_ctrl.temp_ctr\[8\] a_6240_12711# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6068 ts.ts_core.dac_vout_ana_ net14 a_16293_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6069 VPWR res2_n a_6559_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6070 VPWR clknet_0_clk a_7838_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6071 a_9771_18236# a_9576_18267# a_10081_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X6072 a_6658_10966# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X6073 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6074 a_4975_12925# a_4351_12559# a_4867_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6075 a_16609_6575# _061_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6076 _100_ _095_ a_16209_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X6077 a_6447_11837# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6078 ts.ts_core.dac_vout_ana_ net14 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6079 VGND a_6240_12711# _210_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X6080 _098_ a_11606_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X6081 a_4986_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6082 VGND a_13611_4917# net68 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6083 a_10313_2767# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6084 uo_out[6] a_9800_13423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6085 a_9716_13423# ts.o_res\[6\] a_9800_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6086 ts.o_res\[9\] a_12875_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6087 net12 a_18847_16341# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6088 a_4349_17429# a_4131_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6089 a_10313_3855# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6090 ts.ts_ctrl.state\[1\] a_13059_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6091 a_16591_1135# a_16403_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6092 _185_ _177_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6093 VGND net70 a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6094 res1_n a_2439_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6095 _093_ a_10977_9955# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X6096 VPWR a_3111_6794# _024_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6097 a_4126_8983# ts.ts_ctrl.temp_ctr\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6098 a_4513_13621# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6099 a_8448_15975# ts.ts_ctrl.temp_ctr\[15\] a_8590_16150# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X6100 VGND clknet_0_clk a_7838_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6101 a_6690_16911# _185_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
R53 VGND net38 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6102 a_2659_10357# ts.ts_ctrl.temp_ctr\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6103 a_14545_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6104 a_10081_17999# a_9702_18365# a_10009_17999# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X6105 a_11913_16885# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6107 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15952_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6108 a_13967_12711# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.141 ps=1.33 w=0.42 l=0.15
X6109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6110 VPWR a_18234_10927# net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6111 a_17029_2767# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6112 uo_out[4] a_9340_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6113 VPWR _047_ a_9169_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X6114 VPWR ts.ts_ctrl.temp_ctr\[11\] a_6427_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X6115 VPWR _071_ a_10516_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X6116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6117 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6118 a_17673_15599# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6119 a_13326_5719# _140_ a_13463_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6120 VPWR a_5232_6005# _199_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X6121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6122 a_8289_2223# a_7755_2229# a_8194_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6123 _102_ a_11895_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6124 net14 a_17783_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6125 VGND net67 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6126 ts.o_res\[7\] a_7079_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6127 a_11808_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6128 a_17695_8751# a_17507_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6129 a_7815_4917# _153_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X6130 a_7285_12335# ts.ts_ctrl.temp_ctr\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6131 a_14172_3689# a_13091_3317# a_13825_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6132 a_14107_4117# a_13919_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6134 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6135 a_17497_3311# _150_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6136 a_7286_9839# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X6137 a_9169_11721# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X6138 a_9129_15657# a_7939_15285# a_9020_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6139 VPWR a_16863_14735# a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6140 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6141 a_14195_9295# _134_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6142 a_3767_12393# a_3321_12021# a_3671_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6143 a_16315_5487# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6144 VPWR a_14571_11623# a_13836_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6145 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6146 a_11573_7663# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6147 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6148 a_9169_11721# ts.o_res\[12\] a_9340_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6149 a_15951_2919# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6150 VGND clknet_2_2__leaf_clk a_4259_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6151 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6152 VPWR a_1589_10901# a_1479_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6153 _165_ _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6154 a_7759_1135# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6155 a_11101_11721# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X6156 _137_ a_6059_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6157 a_16131_6293# a_15943_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6158 VPWR _059_ _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6159 a_17603_9839# a_17415_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6160 a_14843_13621# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X6161 VGND _187_ a_5905_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6162 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16753_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6163 a_4055_5309# a_3431_4943# a_3947_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6164 VGND _144_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6165 a_15212_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R54 VGND tt_um_hpretl_tt06_tempsens_51.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6166 a_6817_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6167 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12819_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6168 a_6825_13647# ts.ts_ctrl.temp_ctr\[12\] a_6719_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X6169 VPWR a_1551_6807# _009_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X6170 VPWR _164_ _169_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6171 a_1459_14423# _175_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6172 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6174 VGND a_11975_5461# net15 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6175 a_4411_12319# a_4236_12393# a_4590_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6176 a_5423_4917# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X6177 VGND _070_ a_11343_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6178 a_6153_14511# _177_ _190_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6179 VPWR a_16955_4943# a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6181 a_1777_13103# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6182 ts.o_res\[16\] a_7263_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6183 ts.ts_core.dac_vout_ana_ net72 a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6184 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6185 _070_ a_12157_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.247 ps=2.06 w=0.65 l=0.15
X6186 a_8774_16733# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X6187 VGND net67 a_16569_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6188 VGND _087_ a_11696_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
X6189 a_16771_10159# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
X6190 a_2401_5493# a_2235_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6191 a_17029_14735# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6192 ts.ts_core.dac_vout_ana_ net14 a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X6193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6195 a_13832_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6196 VGND a_11207_7637# uio_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6197 _040_ a_10975_17455# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6198 a_5361_6281# _194_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X6199 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6200 a_9573_17999# a_9095_17973# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X6201 VGND net67 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6202 ts.ts_core.dac_vout_ana_ net72 a_9415_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6203 VPWR a_15575_3855# a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6204 VPWR _087_ a_9669_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6205 VPWR a_7937_17429# a_7827_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6206 a_7442_9295# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6207 ts.ts_core.dac_vout_ana_ net72 a_14913_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6208 ts.ts_core.dac_vout_ana_ net15 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6209 VGND net68 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6210 VGND clknet_2_0__leaf_clk a_855_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6211 VPWR a_12127_7093# uio_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6212 VGND a_5043_11636# _031_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6213 VGND net19 a_9913_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6214 a_13928_5487# a_14663_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X6215 a_14882_7983# net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6216 ts.o_res\[19\] a_7539_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6217 a_17143_5205# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6218 VGND _168_ a_3063_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X6219 a_6247_17429# ts.ts_ctrl.temp_ctr\[11\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6220 VGND a_12587_15988# _037_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6221 VPWR a_4279_4123# a_4195_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6222 VPWR a_14287_6031# a_14475_6293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6223 a_10012_15511# ts.o_res\[14\] a_10154_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6224 a_16661_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6225 net53 clknet_2_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6226 a_12319_4777# a_11969_4405# a_12224_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6227 VGND ts.ts_ctrl.state\[2\] a_15229_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6228 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6229 a_15019_9955# a_14986_9849# a_14937_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X6230 a_14374_13799# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X6231 a_13275_6281# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd a_12777_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X6232 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_11803_1679# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6233 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6234 a_12587_15988# _213_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6235 VPWR ts.ts_ctrl.state\[2\] _062_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6236 VPWR a_7539_3829# a_7526_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6237 VGND net69 a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6238 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6239 VPWR a_17699_13799# a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6240 a_11518_8457# _123_ a_11435_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X6241 a_9585_9545# _088_ a_9669_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6242 a_18847_16341# uio_in[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6243 a_8441_5853# a_8397_5461# a_8275_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6244 net16 a_5423_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6245 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6246 ts.ts_core.dac_vout_ana_ net15 a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6248 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd _061_ a_17862_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.175 ps=1.35 w=1 l=0.15
X6249 _008_ _159_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6250 a_11241_13103# _081_ a_11325_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6251 VGND net67 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6253 ts.o_res\[5\] a_7815_13407# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6254 a_11372_11247# ts.o_res\[9\] a_11456_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6255 a_5416_14735# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6256 a_11114_16189# a_10037_15823# a_10952_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6257 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6258 ts.ts_core.dac_vout_ana_ net14 a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6259 a_16683_12015# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6260 ts.ts_core.dac_vout_ana_ net71 a_10335_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6261 a_12157_13799# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X6262 _155_ a_10523_3427# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6263 a_5989_11471# a_5823_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6264 VPWR a_3889_11989# a_3779_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6265 a_12967_15583# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6266 VGND _061_ a_16771_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6267 a_15649_11471# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6268 VPWR a_17507_4399# a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6269 a_13546_13335# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X6270 VGND a_2111_7093# ts.ts_ctrl.temp_ctr\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6271 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6273 a_4135_11445# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X6274 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6275 a_16131_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6277 a_11812_4105# a_12547_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6278 a_11150_9545# _120_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6279 VGND _143_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6280 a_9232_591# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6281 a_1846_4221# a_1407_3855# a_1761_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6282 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6283 VGND a_12679_10071# _087_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X6284 VPWR a_14747_1679# a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6285 a_11812_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6286 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6287 VPWR a_16863_1679# a_17051_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6288 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6289 VPWR a_15123_2197# a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6290 VGND ts.ts_ctrl.state\[2\] a_12447_5540# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X6291 a_10012_5719# _058_ a_10154_5526# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X6292 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6293 a_18787_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.236 pd=1.38 as=0.176 ps=1.84 w=0.65 l=0.15
X6294 VPWR a_17507_6575# a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6295 a_2751_5865# a_2401_5493# a_2656_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6296 VGND net70 a_16863_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6297 a_8084_5853# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6298 VGND net11 _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6299 VPWR a_15399_12711# a_14664_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X6300 a_16131_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6301 a_5502_10749# a_4425_10383# a_5340_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6303 a_18753_10548# ui_in[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6305 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17581_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6306 a_16131_6293# a_15943_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X6307 a_6520_15645# _021_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6308 a_5511_14735# a_4995_14735# a_5416_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6309 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6311 a_16293_5807# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6312 a_3871_16189# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6313 a_13556_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6314 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9227_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6315 ts.ts_ctrl.temp_ctr\[1\] a_11035_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6316 VGND _092_ a_10977_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6317 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6318 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6319 VGND _143_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6320 a_10961_13799# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X6321 a_6427_13621# ts.ts_ctrl.temp_ctr\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X6322 a_12245_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6323 VGND net19 a_9821_16911# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6324 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6325 uo_out[1] a_11456_11247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6326 VGND _151_ a_13551_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6327 VGND net67 a_16127_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6328 a_12427_4399# a_11803_4405# a_12319_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6329 a_11931_7983# _096_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6330 a_9393_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6331 _052_ a_9063_8534# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X6332 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6333 a_10605_3427# a_10331_3671# a_10523_3427# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6334 VGND _143_ ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6335 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6337 a_6557_7637# a_6339_8041# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6338 a_16661_11247# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6339 a_7929_12015# ts.ts_ctrl.temp_ctr\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6340 ts.o_res\[1\] a_8919_5791# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6341 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6342 a_17581_10159# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6343 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16477_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6344 a_2098_7485# a_1021_7119# a_1936_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6345 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6346 a_17673_15599# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6347 a_12819_2223# a_12631_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6348 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6349 a_6247_5461# ts.ts_ctrl.temp_ctr\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6350 a_14418_9071# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6351 a_11969_1679# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6352 _201_ ts.ts_ctrl.temp_ctr\[17\] a_4702_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.091 ps=0.93 w=0.65 l=0.15
X6353 VGND net69 a_16661_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6354 _215_ a_9339_18582# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X6355 VGND a_12596_5461# _058_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X6356 VGND clknet_2_1__leaf_clk a_8767_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6357 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6358 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15465_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6359 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6360 VPWR a_11456_11247# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6361 a_9306_11247# _048_ a_8836_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6362 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6363 a_17191_11445# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X6364 a_10321_9545# _088_ a_10405_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6365 ts.ts_core.o_tempdelay a_10443_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6366 a_13923_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6367 a_13326_5719# net4 a_13540_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6368 a_10513_6273# a_10295_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6369 _159_ a_10294_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X6370 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6372 a_10154_5526# ts.ts_ctrl.temp_ctr\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X6373 a_14567_12015# a_14379_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X6374 a_13601_7983# _113_ a_13183_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6375 a_6339_9129# a_5989_8757# a_6244_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6376 a_16477_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6377 VPWR a_2111_14709# a_2098_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6378 a_1972_3855# a_1573_3855# a_1846_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6380 a_16315_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6381 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6382 VGND a_9061_16665# a_8995_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X6383 VPWR _149_ a_13183_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6384 VPWR net9 a_8449_8790# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X6385 VPWR a_9235_1831# a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6386 a_14292_4719# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6387 a_9287_3829# _153_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X6388 a_4229_6031# ts.ts_ctrl.temp_ctr\[17\] a_4157_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6389 a_15465_13647# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6390 _121_ a_11159_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6391 VGND a_2397_6807# net61 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X6392 a_16793_8751# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6393 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6394 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6395 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6396 VGND clknet_2_2__leaf_clk a_855_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6397 a_14664_12809# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6398 VPWR a_16127_13103# a_16315_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6399 a_9037_13423# ts.ts_ctrl.temp_ctr\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6400 a_6265_15285# a_6099_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6401 a_15487_13909# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6402 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_10313_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6403 VPWR a_7221_7093# a_7251_7446# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6404 a_17673_9071# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6405 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_16293_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6406 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14545_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6407 a_11491_3689# a_11141_3317# a_11396_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6408 a_11969_4405# a_11803_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6409 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6410 VGND _064_ a_14471_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6411 ts.ts_core.capload\[15\].cap.Y net28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6412 a_6339_11471# a_5989_11471# a_6244_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6413 VPWR a_13963_6896# a_13599_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X6414 VGND _094_ _134_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6415 a_7631_17973# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6416 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6417 a_9393_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6418 a_15487_13909# a_15299_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6419 a_17121_14511# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6420 VPWR a_16955_8207# a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6422 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6423 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6424 a_8456_9117# ts.o_res\[19\] a_8235_8790# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6425 ts.ts_core.dac_vout_ana_ net71 a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6426 a_17673_9071# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6427 a_13560_3017# a_14295_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6428 a_14526_3677# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6429 VGND net9 a_13551_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6430 clknet_0_clk a_7286_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6431 a_4588_5807# a_4362_5603# a_4219_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6432 a_16315_13103# a_16127_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X6433 net70 a_17935_13363# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6434 a_2111_11231# a_1936_11305# a_2290_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6435 a_8995_16733# ts.ts_ctrl.temp_ctr\[11\] a_8632_16599# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6436 VGND net72 a_18243_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6437 a_4986_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X6438 a_13633_6353# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6439 a_12797_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6440 VPWR a_10961_13799# _057_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X6441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6442 a_9236_841# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6443 a_14545_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6444 ts.ts_core.dac_vout_ana_ net72 a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6445 a_14384_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R55 tt_um_hpretl_tt06_tempsens_50.LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6446 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6447 a_6557_11713# a_6339_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6448 VGND res1_n a_3177_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6449 ts.ts_core.dac_vout_ana_ net72 a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6450 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6451 VPWR ts.ts_ctrl.temp_ctr\[18\] a_5361_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X6452 VGND net68 a_16863_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6453 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6454 VGND net70 a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6455 a_11808_4943# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6456 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16964_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6457 VPWR ts.ts_ctrl.temp_ctr\[11\] a_5081_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X6458 ts.o_res\[10\] a_12967_15583# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6459 a_8378_3443# a_8695_3553# a_8653_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X6460 a_3299_9269# _163_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X6461 a_6185_2543# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6462 a_17673_9071# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6463 a_7313_4917# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6465 a_16661_12335# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6466 a_18243_7983# _094_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6467 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12797_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6468 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6469 a_6447_8751# a_5823_8757# a_6339_9129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6470 VGND a_10441_15577# a_10375_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X6471 a_12245_1455# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6472 net67 a_17332_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6473 VPWR a_8491_2767# a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6474 VGND a_6427_16341# _021_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6475 VPWR a_2751_15253# a_2493_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.5
X6476 VGND a_5893_5719# net59 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X6477 VGND a_3299_12533# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6478 VGND net54 a_7755_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6479 VPWR a_14295_743# a_13560_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6480 a_14913_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6481 VPWR a_17783_5487# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6482 VPWR net32 ts.ts_core.capload\[4\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6483 a_16311_4943# _140_ a_16465_5193# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6484 a_9214_10159# ts.ts_ctrl.temp_ctr\[3\] a_9128_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X6485 a_10980_2543# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6487 VPWR net4 a_16609_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6488 VGND net67 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6489 VGND a_16180_11989# _067_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6490 a_3321_12021# a_3155_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6491 a_11943_17238# ts.o_res\[13\] a_11484_17063# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X6492 VGND net70 a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6493 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12079_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6494 a_12275_6281# _112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6495 VGND a_18755_3829# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6496 a_4165_5185# a_3947_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6497 VPWR a_16127_2223# a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6498 a_8481_7369# ts.o_res\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6499 VPWR a_1589_7361# a_1479_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6500 VPWR a_17935_13363# net70 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X6501 VGND a_6559_5487# net17 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6502 a_6143_8207# ts.ts_ctrl.temp_ctr\[3\] a_5780_8359# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6503 VGND a_14937_9955# _095_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X6504 a_2375_12247# ts.ts_ctrl.temp_ctr\[4\] a_2609_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6505 a_16863_4719# _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6506 a_9025_13103# ts.ts_ctrl.temp_ctr\[12\] a_8941_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6507 a_6615_15657# a_6099_15285# a_6520_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6508 net55 clknet_2_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6509 _145_ a_8155_4737# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
R56 tt_um_hpretl_tt06_tempsens_46.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6511 VPWR a_12875_14709# a_12862_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6512 VPWR a_16955_7119# a_17143_7381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6513 a_8657_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6514 net15 a_11975_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6515 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6516 a_3859_15823# a_3413_15823# a_3763_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6517 a_9945_6031# a_9779_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6518 VPWR ts.o_res\[8\] a_8217_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6519 VPWR a_12547_743# a_11812_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X6520 ts.ts_core.dac_vout_ana_ net14 a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6521 a_15671_11733# a_15483_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X6522 a_9340_11471# _051_ a_9169_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6523 VPWR a_6945_11225# a_6975_10966# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6524 a_12245_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6525 a_6520_15645# _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6526 a_16187_7895# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6527 a_15304_8207# ts.ts_core.dac.vdac_single.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6528 VPWR a_5729_14977# a_5619_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6529 a_16315_853# a_16127_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6530 VPWR ts.o_res\[10\] a_11101_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6531 VGND clknet_2_3__leaf_clk a_11251_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6532 _133_ a_9597_9955# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X6533 _054_ _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6534 a_13560_841# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6535 a_4680_10383# _031_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6536 VPWR _074_ a_15187_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.5 as=0.0693 ps=0.75 w=0.42 l=0.15
X6537 VPWR a_13735_1135# a_13923_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6539 VPWR ts.ts_ctrl.state\[2\] a_13551_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6540 a_1855_7983# ts.ts_ctrl.temp_ctr\[2\] _160_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X6541 VPWR a_16863_2767# a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6542 VGND net13 a_13905_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X6543 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6544 a_6907_4221# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6545 a_17673_4719# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6546 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6547 a_14101_12559# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.103 ps=1 w=0.42 l=0.15
X6548 ts.ts_core.dac_vout_ana_ net14 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6550 a_11399_1109# ts.ts_core.tempdelay_sync1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6551 a_16170_6895# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6552 a_1479_12925# net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6553 a_9095_17973# a_9298_18251# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X6554 a_3781_17461# a_3615_17461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6556 a_2290_14735# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6557 VPWR a_15943_4943# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6558 a_8022_6575# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6559 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17143_8469# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6560 VGND a_1367_10357# _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6561 a_9687_8751# _089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X6562 a_14189_12559# net11 a_14101_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X6563 a_4126_8983# ts.ts_ctrl.temp_ctr\[16\] a_4446_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6565 _106_ a_8491_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6566 ts.ts_ctrl.temp_ctr\[14\] a_7355_15583# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6567 VPWR a_13086_11159# _078_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X6568 VPWR a_4871_17759# a_4858_17455# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6569 ts.ts_core.dac_vout_ana_ net14 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6570 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_8496_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6571 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6572 VGND _068_ _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6573 a_13560_3017# a_14295_2919# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X6574 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X6575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X6576 a_18763_7271# _139_ a_18937_7147# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6577 a_9781_7369# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6578 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13832_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6579 ts.o_res\[3\] a_7079_9055# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6580 VGND a_3583_14495# a_3517_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6581 VGND ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6582 VGND _074_ _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X6583 a_4512_4943# a_3597_4943# a_4165_5185# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6584 VPWR _095_ a_18243_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6585 a_8573_7983# ts.ts_ctrl.temp_ctr\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6586 a_9415_2223# a_9227_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6588 a_18325_6281# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd _111_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6589 VGND _070_ a_12493_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6590 a_17029_2767# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6591 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6592 _148_ a_17753_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.373 ps=1.75 w=1 l=0.15
X6593 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6594 _150_ a_17017_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6595 VPWR _103_ a_12603_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X6596 a_11053_5719# _058_ a_11216_5603# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6597 a_2695_11721# _164_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X6598 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _061_ a_16793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6599 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_13551_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6600 a_1479_10927# a_855_10933# a_1371_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6601 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6602 VGND ts.o_res\[11\] a_8856_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X6603 VGND a_2111_14709# a_2045_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6604 VPWR _114_ a_13599_6807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X6605 a_11058_9545# _127_ a_10975_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X6606 VGND a_18109_10548# ts.ts_core.dac.vdac_single.en_pupd VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6607 a_9374_15645# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6608 a_10335_3029# net71 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6609 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6610 ts.ts_core.dac_vout_ana_ net14 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6611 a_18763_9447# _139_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6612 a_3045_10933# a_2879_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6613 VGND net67 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6614 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_9393_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6615 a_9414_3311# a_8695_3553# a_8851_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6616 a_10295_6031# a_9945_6031# a_10200_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6617 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6618 a_16661_12335# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6619 a_5541_12559# a_4351_12559# a_5432_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6620 a_16661_11247# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6621 a_16964_13897# a_17699_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6622 VPWR a_5140_15253# _022_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X6623 res2_n a_4279_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6624 VPWR ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16587_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6625 ts.ts_core.dac_vout_ana_ net14 a_11808_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6626 a_10313_3855# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6627 a_10335_1941# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6628 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_13735_1135# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6629 a_11456_11247# ts.o_res\[9\] a_11372_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6630 a_10975_8864# _089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6631 a_9771_18236# a_9615_18141# a_9916_18365# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X6632 a_14475_5205# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X6634 a_15671_11733# a_15483_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6635 VPWR clknet_0_clk a_4986_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6636 net68 a_13611_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6637 _063_ ts.ts_ctrl.state\[0\] a_11601_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X6638 a_14024_8207# a_13643_8207# _140_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6639 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16683_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6640 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17051_14997# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6641 a_4993_10625# a_4775_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6642 VPWR _159_ a_2787_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X6643 VGND _101_ a_12321_12705# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X6644 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6645 VPWR a_16127_2223# a_16315_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6646 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_14453_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6647 a_17029_2767# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6648 VGND _069_ a_11589_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6649 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_11808_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6650 ts.ts_core.dac_vout_ana_ net15 a_7759_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6651 a_14935_1941# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6652 VPWR a_12547_5095# a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6653 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6654 VGND a_3111_6794# _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6655 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6656 VGND a_4513_13621# clknet_2_2__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6657 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6658 a_9100_4765# ts.o_res\[0\] a_8879_4438# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6659 VPWR a_3491_5791# ts.ts_ctrl.temp_ctr\[17\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6660 VGND a_15451_14423# _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X6661 VGND net18 a_3933_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6662 a_12547_4007# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6663 VPWR _157_ _007_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6665 VPWR a_8816_6183# _203_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6666 a_10147_9839# _069_ a_10229_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6667 a_5425_13469# ts.ts_ctrl.temp_ctr\[9\] a_5353_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6668 VPWR a_8468_10357# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6669 a_17121_4943# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6670 VGND a_10012_15511# _217_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X6671 VPWR a_6791_3530# _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6672 net14 a_17783_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6673 a_1761_3855# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6674 VPWR a_10018_4373# a_9945_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6675 a_17051_14997# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6676 a_17051_1941# net15 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6677 VPWR net29 ts.ts_core.capload\[1\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6678 a_6817_591# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6680 VPWR _112_ _114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6681 VGND a_3491_5791# a_3425_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6682 a_9179_6031# ts.ts_ctrl.temp_ctr\[1\] a_8816_6183# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6683 ts.ts_core.dac_vout_ana_ net15 a_17051_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6684 VPWR a_3663_15511# _180_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6685 a_8397_5461# a_8179_5865# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6686 a_4682_8207# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6687 VPWR clknet_2_1__leaf_clk a_6007_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6688 VGND clknet_2_1__leaf_clk a_11803_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6689 a_14663_5461# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6690 a_8958_6031# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X6691 a_6817_591# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6692 a_7313_6005# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6693 uio_out[4] a_11207_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6694 a_14334_3311# a_13257_3317# a_14172_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6695 ts.ts_core.dac_vout_ana_ net14 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6696 a_10335_4117# a_10147_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6697 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6698 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6699 VPWR clknet_2_0__leaf_clk a_855_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6700 _058_ a_12596_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X6701 a_10403_6397# a_9779_6031# a_10295_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6702 VPWR a_3981_16065# a_3871_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6703 VPWR _064_ _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6704 a_16683_10927# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6705 VPWR a_7838_14191# clknet_2_3__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6706 a_18763_8359# _150_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6707 a_16569_1455# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6708 a_3779_12015# a_3155_12021# a_3671_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6709 net20 a_4680_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6710 VPWR a_1367_10357# _011_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X6711 VGND net69 a_16495_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6712 a_16477_12559# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6713 VPWR _087_ a_9045_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6714 a_16960_13647# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6715 VGND net70 a_17673_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6716 a_13238_4765# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6717 a_15321_7663# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6718 a_16293_13423# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6719 a_17581_10159# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6720 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6721 a_14475_6293# a_14287_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6722 _191_ a_5271_13216# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6723 a_9284_8207# ts.o_res\[17\] a_9063_8534# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6724 a_7749_13481# a_6559_13109# a_7640_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6725 VGND a_11975_5461# net15 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6726 a_14660_12559# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6727 a_7293_13077# a_7075_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6728 a_12135_14735# a_11619_14735# a_12040_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6729 a_12596_5461# a_12447_5540# a_12892_5603# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6730 VPWR _075_ a_8481_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6731 a_15125_10383# _073_ a_14857_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X6732 a_6829_1455# ts.ts_core.dcdel_capnode_ana_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6733 a_4036_17821# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6734 a_6769_17821# _177_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6735 VGND _112_ a_12591_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6737 a_13257_3317# a_13091_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6738 VGND net68 a_11808_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6739 a_13546_10535# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X6740 VPWR _114_ a_6690_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X6741 ts.o_res\[14\] a_11127_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6742 ts.ts_core.dac_vout_ana_ net72 a_10980_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6743 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6744 a_15304_8207# net47 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6745 a_16775_7663# a_16587_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X6746 a_8413_3677# a_8378_3443# a_8175_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X6747 a_8836_10901# ts.o_res\[0\] a_9658_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6748 a_9089_3677# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X6749 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6750 a_6631_4399# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6751 VPWR net70 a_16127_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6752 VPWR net10 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6753 VGND net17 a_9545_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6754 VGND _084_ a_12149_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X6755 a_14195_9295# _133_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6756 a_18755_3829# _142_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X6757 a_16212_4719# ts.ts_ctrl.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6758 VGND _121_ a_12079_8457# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X6759 VGND clknet_2_2__leaf_clk a_6007_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6760 a_3503_10927# a_2879_10933# a_3395_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6761 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_17121_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6762 a_15948_9295# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6764 a_2098_15101# a_1021_14735# a_1936_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6765 _094_ a_15535_10357# a_15315_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6766 a_6427_13621# ts.ts_ctrl.temp_ctr\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X6767 a_10012_5719# _112_ a_10154_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6768 VGND net67 a_16109_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6769 a_10055_10927# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X6770 VGND net67 a_11969_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6771 net69 a_18234_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6772 ts.ts_core.dac_vout_ana_ net15 a_17029_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6773 a_7394_12886# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X6774 a_7737_1455# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6775 VPWR a_8448_4007# _222_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6776 VPWR a_14347_3615# ts.ts_ctrl.state\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6777 a_13928_5487# a_14663_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6778 a_16315_13103# a_16127_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6779 a_4055_5309# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6780 VGND a_13599_6807# _115_ VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6781 _092_ a_9503_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X6782 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15487_13909# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6783 a_9188_4943# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6784 a_7775_8534# ts.o_res\[18\] a_7703_8534# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6785 a_6339_11471# a_5823_11471# a_6244_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6786 VGND _069_ a_11129_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6787 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6788 VPWR _065_ ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X6789 ts.o_res\[4\] a_5515_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6790 a_9501_5185# a_9283_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6791 VPWR ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd a_16955_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6792 a_2305_10535# a_2401_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.5
X6793 a_14828_14557# a_14379_14191# a_14526_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6794 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6795 a_7247_4943# ts.ts_ctrl.temp_ctr\[18\] a_6884_5095# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6796 VPWR a_6427_13621# _187_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X6797 VPWR a_16495_10927# a_16683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6798 a_9500_12015# ts.o_res\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6799 VGND net70 a_17121_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6800 a_1479_8751# a_855_8757# a_1371_9129# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6801 a_7394_12559# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X6802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6803 a_9585_9545# _091_ a_9503_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6804 _051_ net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6805 VPWR a_16955_4943# a_17143_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6806 a_7313_4917# _211_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6807 a_4683_13077# ts.ts_ctrl.temp_ctr\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6808 a_17695_15279# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6809 a_7775_8207# a_7521_8534# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X6810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6811 ts.ts_core.tempdelay_async ts.ts_core.dcdel_out_n VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6812 VPWR a_8919_5791# a_8906_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6813 net8 a_8399_18543# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X6814 ts.ts_core.dac_vout_ana_ net14 a_15308_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6815 VPWR a_18763_8359# _151_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X6816 clknet_2_2__leaf_clk a_4513_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6817 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_17121_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6818 a_10334_18365# a_9615_18141# a_9771_18236# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6819 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_9232_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6820 VPWR a_5423_4917# net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6821 clknet_2_0__leaf_clk a_4986_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6822 a_12181_7663# _093_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6823 a_9339_18909# a_9085_18582# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X6824 VPWR clknet_2_3__leaf_clk a_7203_17461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6825 VPWR a_17507_4399# a_17695_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6826 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6827 a_10952_15823# a_10037_15823# a_10605_16065# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6828 uio_out[7] a_14717_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6829 VPWR a_17191_11445# _074_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6830 a_16683_10927# a_16495_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6831 a_17121_14511# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6832 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_13556_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6833 VGND net68 a_17673_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6834 a_13963_6896# _095_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6835 a_9770_10383# ts.o_res\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X6836 VPWR a_4512_4943# a_4687_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6837 a_16964_13897# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6838 VGND _050_ _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6839 VPWR net20 a_8399_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6840 a_17143_5205# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6841 VGND ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref a_16955_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6842 clknet_2_3__leaf_clk a_7838_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X6843 VPWR ts.ts_ctrl.state\[2\] a_12447_5540# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X6844 net67 a_17332_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6845 clknet_2_1__leaf_clk a_8022_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6846 VGND a_6791_3530# _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6847 a_10313_3855# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6848 VPWR _113_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6849 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd a_17673_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6850 _076_ a_9770_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X6851 VGND net67 a_14379_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6852 a_12127_7093# a_12493_7369# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6853 a_17753_9545# _098_ a_17681_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
X6854 ts.ts_core.dac_vout_ana_ net15 a_13556_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6855 VGND net67 a_14545_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6856 a_12537_4373# a_12319_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6857 a_16315_5487# a_16127_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6858 a_11553_5825# _146_ a_11467_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6859 res2_n a_4279_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6860 a_4972_4777# a_4057_4405# a_4625_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6861 VPWR a_17507_6575# a_17695_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6863 a_7252_12711# ts.ts_ctrl.temp_ctr\[5\] a_7394_12886# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X6864 a_9971_743# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6865 a_12231_3615# a_12056_3689# a_12410_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6866 a_7263_4703# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6868 clknet_2_0__leaf_clk a_4986_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6869 VPWR a_11709_3285# a_11599_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6870 VPWR a_13825_3285# a_13715_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6871 VGND a_18763_7271# _149_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X6872 VGND clknet_2_0__leaf_clk a_5823_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6873 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6874 a_10292_15823# _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6875 VPWR _140_ a_17141_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.117 ps=1.24 w=1 l=0.15
X6876 VGND net67 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6877 a_18753_10548# ui_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6878 a_5432_12559# a_4517_12559# a_5085_12801# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6879 a_15212_2767# ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6880 VPWR _059_ a_12691_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X6881 a_13183_7663# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X6882 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _061_ a_15321_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6883 a_7815_13407# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6884 a_11931_7983# a_11573_7663# a_11207_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6885 a_16354_9071# _065_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6886 a_9393_2543# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6887 VGND net67 a_15304_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6888 a_1021_8757# a_855_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6889 VPWR a_7365_15975# net66 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6890 a_17143_7381# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6891 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6892 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X6893 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6894 a_7258_9117# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6895 VGND _061_ a_13643_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.04 as=0.109 ps=1.36 w=0.42 l=0.15
X6896 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_14296_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6897 a_5094_11293# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X6898 uo_out[2] a_11272_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X6899 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6900 VGND a_18848_13621# net10 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6901 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6902 a_14418_9071# _097_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6903 VGND ts.ts_ctrl.temp_ctr\[5\] _166_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6904 a_11969_1679# net71 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6905 a_4680_10383# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6906 a_7937_17429# a_7719_17833# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6907 a_6645_16367# net66 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6908 a_1936_14735# a_1021_14735# a_1589_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6909 VGND _058_ a_11573_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6910 _068_ a_13603_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6911 VGND net16 a_6785_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6912 VPWR a_15483_11471# a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6913 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15763_4117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6914 VPWR a_8447_6196# _028_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6915 a_2748_14557# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6916 a_3852_4943# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6917 ts.ts_ctrl.temp_ctr\[3\] a_2111_9055# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6918 VGND net18 a_1633_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6919 VPWR ts.ts_core.dcdel_capnode_ana_ ts.ts_core.capload\[3\].cap.Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6920 ts.ts_core.capload\[6\].cap.Y net34 a_6461_591# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6921 a_11851_12247# ts.o_res\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6922 a_11435_8207# _122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X6923 a_10984_2223# a_11719_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6924 VPWR a_11803_1679# a_11991_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6925 a_3668_8207# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6926 a_11672_17821# _040_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6927 a_16945_4399# ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6928 _112_ ts.ts_ctrl.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6929 a_6033_13469# _187_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6930 VPWR ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_12631_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6931 a_16315_2223# net72 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6932 a_1589_12801# a_1371_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6933 a_12445_15253# a_12227_15657# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6934 VGND clknet_2_2__leaf_clk a_3615_17461# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6935 a_6563_16687# _186_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X6936 VPWR a_9235_1831# a_8500_1929# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X6937 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_13919_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6938 a_10607_12809# _088_ a_10689_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6939 ts.ts_core.dac_vout_ana_ net15 a_11812_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6940 a_3435_12559# _167_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X6941 VGND ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_14085_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X6944 a_4858_17455# a_3781_17461# a_4696_17833# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6945 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_15483_1135# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6946 a_16683_10927# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6947 a_3307_13799# ts.ts_ctrl.temp_ctr\[8\] a_3481_13675# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6948 _174_ _172_ a_3329_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X6949 a_5232_6005# ts.ts_ctrl.temp_ctr\[17\] a_5455_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X6950 _141_ a_16465_5193# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6951 a_17673_9071# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6952 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6953 _129_ a_7203_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6954 VGND ts.ts_ctrl.temp_ctr\[10\] a_5425_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6955 a_8632_16599# ts.o_res\[11\] a_8774_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6956 VPWR a_6792_7271# _204_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6957 _143_ _122_ a_13183_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6958 a_16569_10383# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6959 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6960 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6961 a_12313_12234# _084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6962 VPWR a_12079_1135# a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X6963 a_9393_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6964 VPWR net3 a_16793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6965 a_17332_3829# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6966 VGND a_4986_7119# clknet_2_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6967 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_9236_841# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6968 a_14660_12559# net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X6969 a_14664_12809# a_15399_12711# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6970 a_14913_1679# net72 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6971 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref a_10147_1679# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6972 VPWR clknet_2_3__leaf_clk a_7939_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6973 a_15123_2197# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6974 VPWR clknet_2_0__leaf_clk a_3247_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6975 a_7183_13103# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6977 VGND net67 a_7737_1455# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X6978 ts.ts_core.dac_vout_ana_ net71 a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6979 VPWR a_18335_2223# net72 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6980 a_14107_4117# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6981 VPWR net10 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6982 VPWR _177_ a_6883_14887# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X6983 ts.ts_core.dac_vout_ana_ net15 a_6817_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6984 a_14418_9071# _108_ a_14584_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6985 a_9889_13621# _154_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6986 VPWR a_14747_1679# a_14935_1941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X6987 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16569_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6988 VGND a_18756_15797# net11 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6989 VGND net69 a_16661_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6990 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd _065_ a_14882_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X6991 a_16180_11989# net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X6992 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X6993 a_11808_4943# net15 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6994 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6995 a_16131_6293# net14 ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6996 VPWR a_4986_7119# clknet_2_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6997 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd a_16775_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X6998 a_11812_4105# a_12547_4007# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.244 pd=2.4 as=0.127 ps=1.21 w=0.94 l=0.15
X6999 VGND ts.ts_ctrl.state\[0\] a_10523_3427# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7000 VPWR a_7286_9839# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7001 VPWR ts.o_res\[7\] a_9500_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7002 uo_out[7] a_9112_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7003 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7004 a_12896_12559# net9 a_12321_12705# VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X7005 a_9889_13621# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X7006 a_10668_7119# a_10625_7352# a_10596_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X7007 a_10009_17999# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X7008 a_13560_3017# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7009 clknet_2_3__leaf_clk a_7838_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7010 a_17121_8207# ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7011 a_17051_14997# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7012 VPWR net64 a_1762_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X7013 VPWR _065_ _140_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7014 a_8856_10383# net8 a_8468_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7015 VGND clknet_2_1__leaf_clk a_10975_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7016 VGND clknet_2_1__leaf_clk a_13091_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7017 a_4512_4943# a_3431_4943# a_4165_5185# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7018 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7019 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7020 a_14913_1679# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7021 a_17029_1679# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7022 a_7615_12559# ts.ts_ctrl.temp_ctr\[5\] a_7252_12711# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7023 net72 a_18335_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7024 a_5773_14735# a_5729_14977# a_5607_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X7025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7026 a_9232_591# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7027 a_9112_11989# _051_ a_9500_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7029 a_14500_8751# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X7030 VGND net69 a_15649_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7031 a_4328_8207# a_3247_8207# a_3981_8449# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7032 _059_ net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7033 VPWR a_10012_5719# _157_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X7034 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7035 a_5269_15599# _186_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X7036 a_8657_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7037 VGND a_7252_12711# _207_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X7038 _138_ a_5179_16367# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7039 uo_out[3] a_8468_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7040 a_16393_5193# ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7041 a_11969_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7042 a_6975_10966# ts.o_res\[7\] a_6516_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X7043 VPWR a_12332_17833# a_12507_17759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7044 VPWR _066_ a_14177_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X7045 a_3686_4221# a_3247_3855# a_3601_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7046 ts.ts_core.dac_vout_ana_ net14 a_16591_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
R57 VPWR ts.ts_core.capload\[0\].cap_22.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7047 VGND _050_ a_11724_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X7048 a_16683_10927# a_16495_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7049 a_9800_13423# _057_ a_10068_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7050 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7051 a_6557_7637# a_6339_8041# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7052 VPWR a_14287_4943# a_14475_5205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.244 ps=2.4 w=0.94 l=0.15
X7053 ts.o_res\[2\] a_7079_7967# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7054 a_17029_14735# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7055 a_8657_2767# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7056 VGND ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd a_17507_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7058 VPWR a_6669_12533# a_6699_12886# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7059 a_16293_13423# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7060 VPWR a_7263_4703# a_7250_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7061 net17 a_6559_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7062 VGND a_4126_8983# _194_ VGND sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0878 ps=0.92 w=0.65 l=0.15
X7063 a_6447_8751# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7064 ts.ts_core.dac_vout_ana_ net14 a_14567_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7065 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref _144_ a_13845_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7066 a_12245_1455# ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R58 VPWR uio_oe[5] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7067 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd _065_ a_16354_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X7068 a_16293_591# net14 ts.ts_core.dac_vout_ana_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7069 VGND a_14717_9545# uio_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7070 VPWR a_8022_6575# clknet_2_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7071 a_15115_9955# _067_ a_15019_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X7072 a_13059_4703# a_12884_4777# a_13238_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7073 a_9687_10633# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X7074 VGND a_4135_11445# net18 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7075 VGND a_16640_14165# _073_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X7076 a_7442_6941# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7077 a_6185_17161# _182_ a_6101_17161# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7078 VGND net69 a_16960_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7079 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_16293_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7081 VGND a_4219_5461# _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X7082 a_11456_11247# _050_ a_11285_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7083 a_3613_10901# a_3395_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7084 a_9770_10633# _075_ a_9770_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X7085 VPWR a_12079_1135# a_12267_1135# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7086 a_8877_9269# _211_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X7087 a_9415_2223# a_9227_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.33 as=0.127 ps=1.21 w=0.94 l=0.15
X7088 VPWR a_15951_2919# a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.16 ps=1.33 w=0.94 l=0.15
X7089 ts.ts_core.dac_vout_ana_ ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd a_13924_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7090 a_9182_15279# a_8105_15285# a_9020_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7091 VPWR _071_ a_10405_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7092 VPWR a_4513_13621# clknet_2_2__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7093 a_10441_5785# ts.ts_ctrl.temp_ctr\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7094 ts.ts_core.dac_vout_ana_ net14 a_14453_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7095 a_14852_8751# _100_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7096 a_6983_15797# ts.ts_ctrl.temp_ctr\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7097 a_8941_13103# _082_ a_9025_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7098 VGND a_6331_12234# _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7099 ts.ts_ctrl.temp_ctr\[2\] a_2111_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X7100 a_9658_11247# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7101 a_11767_17833# a_11251_17461# a_11672_17821# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7102 _131_ a_7847_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7103 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7104 VPWR a_10605_16065# a_10495_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7105 a_5315_11293# ts.ts_ctrl.temp_ctr\[4\] a_4952_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7106 VPWR net69 a_16403_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7108 a_2271_4221# a_1407_3855# a_2014_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7109 ts.ts_ctrl.temp_ctr\[8\] a_3583_14495# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X7110 net69 a_18234_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7111 VPWR ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref a_15575_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7112 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X7113 VPWR a_15951_2919# a_15216_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7114 ts.ts_core.dac_vout_ana_ net72 a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7116 a_12493_7369# _110_ a_12493_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7117 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X7118 ts.ts_core.dac_vout_ana_ net72 a_14388_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7119 a_17695_15279# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7120 a_4799_9071# _172_ _193_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X7121 a_11977_13103# ts.ts_ctrl.temp_ctr\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7122 a_2969_5461# a_2751_5865# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7123 VPWR _068_ a_14707_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X7124 a_10391_14709# a_10216_14735# a_10570_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7125 a_3812_3855# a_3413_3855# a_3686_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7126 VPWR _051_ _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7127 a_14295_743# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7128 ts.ts_core.dac_vout_ana_ net14 a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
X7129 clknet_0_clk a_7286_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7130 a_12537_4373# a_12319_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7131 a_6904_8041# a_5823_7669# a_6557_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7132 VPWR _070_ a_11593_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7133 _113_ a_12275_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X7134 VPWR clknet_2_3__leaf_clk a_9043_16911# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7135 net19 a_8399_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7136 VPWR a_16043_8359# a_15308_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7137 a_11812_5193# a_12547_5095# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7138 VGND a_18234_10927# net69 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7139 a_8919_5791# net17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7140 a_3491_5791# a_3316_5865# a_3670_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7141 a_3871_16189# a_3247_15823# a_3763_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7142 a_6719_13647# ts.ts_ctrl.temp_ctr\[13\] a_6623_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X7143 VGND a_3853_7093# _195_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7144 VPWR _143_ a_17497_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7145 ts.ts_ctrl.temp_ctr\[17\] a_3491_5791# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X7146 a_16043_7271# net67 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7147 a_2778_11471# _168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X7148 ts.ts_core.dac_vout_ana_ net14 a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.33 w=1 l=0.15
R59 VGND tt_um_hpretl_tt06_tempsens_48.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7149 a_5594_12925# a_4517_12559# a_5432_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7150 a_8175_3285# a_8378_3443# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X7151 a_9415_1135# ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7152 a_12335_15279# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7153 a_14296_4399# a_15031_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7154 _211_ a_7815_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X7155 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_15671_11733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7156 a_13825_3285# a_13607_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7157 ts.ts_core.dac_vout_ana_ ts.ts_core.dac_vout_ana_ a_17695_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7158 _156_ _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7159 a_18774_3311# a_18597_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7160 VPWR a_17783_5487# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7161 VPWR a_11803_2767# a_11991_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7162 a_17673_9071# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X7163 VGND a_4952_11159# _206_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X7164 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_10313_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7165 a_12570_12809# _102_ a_12321_12705# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7166 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref _141_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7167 _164_ a_3299_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7168 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7169 net67 a_17332_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.113 ps=1.38 w=0.42 l=0.15
X7170 VGND clknet_2_3__leaf_clk a_11619_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7171 a_16640_14165# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X7172 VPWR a_8491_2767# a_8679_3029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.21 as=0.127 ps=1.21 w=0.94 l=0.15
X7173 a_7838_14191# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X7174 a_17017_4399# net2 a_16863_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X7176 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7177 VGND ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd a_16293_2543# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 uio_in[7] VGND 0.182f
C1 uio_in[6] VGND 0.182f
C2 uio_in[5] VGND 0.182f
C3 uio_in[4] VGND 0.182f
C4 ena VGND 0.182f
C5 uio_oe[3] VGND 1.49f
C6 uio_oe[6] VGND 0.888f
C7 uio_oe[5] VGND 1.75f
C8 uio_oe[1] VGND 0.917f
C9 uio_out[1] VGND 1.66f
C10 uio_out[0] VGND 1.3f
C11 uio_oe[0] VGND 1.21f
C12 ui_in[4] VGND 2.74f
C13 ui_in[5] VGND 3f
C14 ui_in[2] VGND 2.56f
C15 ui_in[3] VGND 1.99f
C16 rst_n VGND 1.06f
C17 uio_out[6] VGND 3.55f
C18 uio_out[4] VGND 3.77f
C19 uio_out[5] VGND 2.86f
C20 uio_out[7] VGND 2.94f
C21 clk VGND 7.07f
C22 ui_in[1] VGND 1.62f
C23 uo_out[3] VGND 4.5f
C24 uo_out[1] VGND 4.21f
C25 uo_out[0] VGND 4.26f
C26 uo_out[2] VGND 4.07f
C27 uo_out[4] VGND 4.45f
C28 ui_in[0] VGND 2.56f
C29 uo_out[7] VGND 3.75f
C30 uo_out[5] VGND 3.48f
C31 uo_out[6] VGND 3.37f
C32 uio_in[0] VGND 1.24f
C33 ui_in[7] VGND 1.76f
C34 uio_in[3] VGND 1.45f
C35 uio_in[1] VGND 1.33f
C36 uio_in[2] VGND 1.8f
C37 uio_out[2] VGND 1.09f
C38 uio_oe[2] VGND 1.09f
C39 uio_out[3] VGND 1.09f
C40 ui_in[6] VGND 1.15f
C41 uio_oe[7] VGND 0.972f
C42 uio_oe[4] VGND 1.09f
C43 VPWR VGND 1.34p
C44 tt_um_hpretl_tt06_tempsens_42.HI VGND 0.415f $ **FLOATING
C45 tt_um_hpretl_tt06_tempsens_50.LO VGND 0.479f $ **FLOATING
C46 tt_um_hpretl_tt06_tempsens_49.LO VGND 0.479f $ **FLOATING
C47 a_16293_591# VGND 0.824f $ **FLOATING
C48 a_13556_591# VGND 0.824f $ **FLOATING
C49 a_11808_591# VGND 0.824f $ **FLOATING
C50 a_16315_853# VGND 1.18f $ **FLOATING
C51 a_13560_841# VGND 1.18f $ **FLOATING
C52 a_9232_591# VGND 0.824f $ **FLOATING
C53 a_11812_841# VGND 1.18f $ **FLOATING
C54 ts.ts_core.capload\[11\].cap.Y VGND 0.281f $ **FLOATING
C55 ts.ts_core.capload\[1\].cap_29.HI VGND 0.415f $ **FLOATING
C56 a_9236_841# VGND 1.18f $ **FLOATING
C57 ts.ts_core.capload\[5\].cap.Y VGND 0.281f $ **FLOATING
C58 a_16127_591# VGND 1.46f $ **FLOATING
C59 a_14295_743# VGND 1.46f $ **FLOATING
C60 a_12547_743# VGND 1.46f $ **FLOATING
C61 a_9971_743# VGND 1.46f $ **FLOATING
C62 ts.ts_core.capload\[4\].cap_32.HI VGND 0.415f $ **FLOATING
C63 a_6817_591# VGND 0.824f $ **FLOATING
C64 a_6839_853# VGND 1.18f $ **FLOATING
C65 ts.ts_core.capload\[6\].cap.Y VGND 0.281f $ **FLOATING
C66 ts.ts_core.capload\[15\].cap.Y VGND 0.281f $ **FLOATING
C67 ts.ts_core.capload\[0\].cap.Y VGND 0.281f $ **FLOATING
C68 tt_um_hpretl_tt06_tempsens_40.HI VGND 0.415f $ **FLOATING
C69 a_6651_591# VGND 1.46f $ **FLOATING
C70 a_16591_1135# VGND 1.18f $ **FLOATING
C71 a_13923_1135# VGND 1.18f $ **FLOATING
C72 tt_um_hpretl_tt06_tempsens_44.HI VGND 0.415f $ **FLOATING
C73 a_16569_1455# VGND 0.824f $ **FLOATING
C74 a_12267_1135# VGND 1.18f $ **FLOATING
C75 a_16403_1135# VGND 1.46f $ **FLOATING
C76 a_13901_1455# VGND 0.824f $ **FLOATING
C77 a_13735_1135# VGND 1.46f $ **FLOATING
C78 a_12245_1455# VGND 0.824f $ **FLOATING
C79 a_12079_1135# VGND 1.46f $ **FLOATING
C80 a_9415_1135# VGND 1.18f $ **FLOATING
C81 a_7759_1135# VGND 1.18f $ **FLOATING
C82 net28 VGND 1.06f $ **FLOATING
C83 ts.ts_core.capload\[8\].cap.Y VGND 0.281f $ **FLOATING
C84 a_9393_1455# VGND 0.824f $ **FLOATING
C85 a_9227_1135# VGND 1.46f $ **FLOATING
C86 a_7737_1455# VGND 0.824f $ **FLOATING
C87 a_7571_1135# VGND 1.46f $ **FLOATING
C88 ts.ts_core.capload\[10\].cap.Y VGND 0.281f $ **FLOATING
C89 ts.ts_core.capload\[4\].cap.Y VGND 0.281f $ **FLOATING
C90 ts.ts_core.capload\[1\].cap.Y VGND 0.281f $ **FLOATING
C91 ts.ts_core.capload\[14\].cap.Y VGND 0.281f $ **FLOATING
C92 ts.ts_core.capload\[9\].cap.Y VGND 0.281f $ **FLOATING
C93 a_18243_1135# VGND 0.988f $ **FLOATING
C94 a_15483_1135# VGND 0.988f $ **FLOATING
C95 a_11399_1109# VGND 0.788f $ **FLOATING
C96 a_11141_1109# VGND 0.794f $ **FLOATING
C97 a_11045_1367# VGND 0.553f $ **FLOATING
C98 net32 VGND 1.56f $ **FLOATING
C99 net29 VGND 1.82f $ **FLOATING
C100 ts.ts_core.capload\[15\].cap_28.HI VGND 0.415f $ **FLOATING
C101 ts.ts_core.capload\[3\].cap.Y VGND 0.281f $ **FLOATING
C102 tt_um_hpretl_tt06_tempsens_43.HI VGND 0.415f $ **FLOATING
C103 a_17029_1679# VGND 0.824f $ **FLOATING
C104 a_14913_1679# VGND 0.824f $ **FLOATING
C105 a_17051_1941# VGND 1.18f $ **FLOATING
C106 a_11969_1679# VGND 0.824f $ **FLOATING
C107 a_10313_1679# VGND 0.824f $ **FLOATING
C108 a_8496_1679# VGND 0.824f $ **FLOATING
C109 a_14935_1941# VGND 1.18f $ **FLOATING
C110 a_11991_1941# VGND 1.18f $ **FLOATING
C111 a_10335_1941# VGND 1.18f $ **FLOATING
C112 a_8500_1929# VGND 1.18f $ **FLOATING
C113 a_16863_1679# VGND 1.46f $ **FLOATING
C114 a_14747_1679# VGND 1.46f $ **FLOATING
C115 a_13643_1679# VGND 0.525f $ **FLOATING
C116 a_11803_1679# VGND 1.46f $ **FLOATING
C117 a_10147_1679# VGND 1.46f $ **FLOATING
C118 a_9235_1831# VGND 1.46f $ **FLOATING
C119 net36 VGND 2.68f $ **FLOATING
C120 ts.ts_core.capload\[8\].cap_36.HI VGND 0.415f $ **FLOATING
C121 ts.ts_core.capload\[10\].cap_23.HI VGND 0.415f $ **FLOATING
C122 net23 VGND 1.09f $ **FLOATING
C123 net33 VGND 1.98f $ **FLOATING
C124 ts.ts_core.capload\[5\].cap_33.HI VGND 0.415f $ **FLOATING
C125 net24 VGND 3.08f $ **FLOATING
C126 ts.ts_core.capload\[11\].cap_24.HI VGND 0.415f $ **FLOATING
C127 ts.ts_core.capload\[3\].cap_31.HI VGND 0.415f $ **FLOATING
C128 ts.ts_core.capload\[13\].cap.Y VGND 0.281f $ **FLOATING
C129 ts.ts_core.dcdel_out_n VGND 0.794f $ **FLOATING
C130 net31 VGND 1.24f $ **FLOATING
C131 net22 VGND 1.35f $ **FLOATING
C132 ts.ts_core.capload\[0\].cap_22.HI VGND 0.415f $ **FLOATING
C133 tt_um_hpretl_tt06_tempsens_39.HI VGND 0.415f $ **FLOATING
C134 a_16315_2223# VGND 1.18f $ **FLOATING
C135 a_14388_2223# VGND 1.18f $ **FLOATING
C136 a_12819_2223# VGND 1.18f $ **FLOATING
C137 a_10984_2223# VGND 1.18f $ **FLOATING
C138 a_9415_2223# VGND 1.18f $ **FLOATING
C139 a_16293_2543# VGND 0.824f $ **FLOATING
C140 a_16127_2223# VGND 1.46f $ **FLOATING
C141 a_15123_2197# VGND 1.46f $ **FLOATING
C142 a_14384_2543# VGND 0.824f $ **FLOATING
C143 a_12797_2543# VGND 0.824f $ **FLOATING
C144 a_12631_2223# VGND 1.46f $ **FLOATING
C145 a_11719_2197# VGND 1.46f $ **FLOATING
C146 a_10980_2543# VGND 0.824f $ **FLOATING
C147 a_9393_2543# VGND 0.824f $ **FLOATING
C148 a_9227_2223# VGND 1.46f $ **FLOATING
C149 ts.ts_core.tempdelay_sync1 VGND 2.16f $ **FLOATING
C150 a_8109_2223# VGND 0.23f $ **FLOATING
C151 a_18937_2442# VGND 0.524f $ **FLOATING
C152 a_18335_2223# VGND 0.988f $ **FLOATING
C153 net72 VGND 13.1f $ **FLOATING
C154 a_8619_2223# VGND 0.609f $ **FLOATING
C155 a_8787_2197# VGND 0.817f $ **FLOATING
C156 a_8194_2223# VGND 0.626f $ **FLOATING
C157 a_8362_2197# VGND 0.581f $ **FLOATING
C158 a_7921_2229# VGND 1.43f $ **FLOATING
C159 ts.ts_core.tempdelay_async VGND 1.64f $ **FLOATING
C160 a_7755_2229# VGND 1.81f $ **FLOATING
C161 ts.ts_core.capload\[2\].cap_30.HI VGND 0.415f $ **FLOATING
C162 ts.ts_core.capload\[7\].cap_35.HI VGND 0.415f $ **FLOATING
C163 ts.ts_core.capload\[13\].cap_26.HI VGND 0.415f $ **FLOATING
C164 net26 VGND 1.33f $ **FLOATING
C165 ts.ts_core.capload\[12\].cap_25.HI VGND 0.415f $ **FLOATING
C166 net34 VGND 1.47f $ **FLOATING
C167 ts.ts_core.capload\[6\].cap_34.HI VGND 0.415f $ **FLOATING
C168 ts.ts_core.capload\[12\].cap.Y VGND 0.281f $ **FLOATING
C169 ts.ts_core.capload\[2\].cap.Y VGND 0.281f $ **FLOATING
C170 net25 VGND 0.938f $ **FLOATING
C171 net30 VGND 1.44f $ **FLOATING
C172 a_17029_2767# VGND 0.824f $ **FLOATING
C173 a_15212_2767# VGND 0.824f $ **FLOATING
C174 a_13556_2767# VGND 0.824f $ **FLOATING
C175 a_11969_2767# VGND 0.824f $ **FLOATING
C176 a_10313_2767# VGND 0.824f $ **FLOATING
C177 a_8657_2767# VGND 0.824f $ **FLOATING
C178 a_17051_3029# VGND 1.18f $ **FLOATING
C179 a_15216_3017# VGND 1.18f $ **FLOATING
C180 a_13560_3017# VGND 1.18f $ **FLOATING
C181 a_11991_3029# VGND 1.18f $ **FLOATING
C182 a_10335_3029# VGND 1.18f $ **FLOATING
C183 ts.ts_core.capload\[9\].cap_37.HI VGND 0.415f $ **FLOATING
C184 a_8679_3029# VGND 1.18f $ **FLOATING
C185 net54 VGND 1.07f $ **FLOATING
C186 a_18937_2932# VGND 0.524f $ **FLOATING
C187 a_16863_2767# VGND 1.46f $ **FLOATING
C188 a_15951_2919# VGND 1.46f $ **FLOATING
C189 a_14295_2919# VGND 1.46f $ **FLOATING
C190 a_11803_2767# VGND 1.46f $ **FLOATING
C191 a_10147_2767# VGND 1.46f $ **FLOATING
C192 a_8491_2767# VGND 1.46f $ **FLOATING
C193 net37 VGND 2.02f $ **FLOATING
C194 ts.ts_core.capload\[14\].cap_27.HI VGND 0.415f $ **FLOATING
C195 net27 VGND 1.77f $ **FLOATING
C196 ts.ts_core.capload\[7\].cap.Y VGND 0.281f $ **FLOATING
C197 net35 VGND 1.15f $ **FLOATING
C198 ts.ts_core.dcdel_capnode_ana_ VGND 12.2f $ **FLOATING
C199 a_19057_3311# VGND 0.227f $ **FLOATING
C200 a_18880_3311# VGND 0.498f $ **FLOATING
C201 a_18774_3311# VGND 0.578f $ **FLOATING
C202 a_18597_3311# VGND 0.5f $ **FLOATING
C203 a_18278_3311# VGND 0.535f $ **FLOATING
C204 a_13715_3311# VGND 0.168f $ **FLOATING
C205 a_13512_3677# VGND 0.259f $ **FLOATING
C206 a_11599_3311# VGND 0.168f $ **FLOATING
C207 a_8996_3311# VGND 0.168f $ **FLOATING
C208 a_11396_3677# VGND 0.259f $ **FLOATING
C209 a_15571_3311# VGND 0.553f $ **FLOATING
C210 a_15465_3311# VGND 0.794f $ **FLOATING
C211 a_15229_3311# VGND 0.788f $ **FLOATING
C212 a_14172_3689# VGND 0.736f $ **FLOATING
C213 a_14347_3615# VGND 1.54f $ **FLOATING
C214 a_13607_3689# VGND 0.714f $ **FLOATING
C215 a_13825_3285# VGND 0.653f $ **FLOATING
C216 a_13257_3317# VGND 1.57f $ **FLOATING
C217 a_13091_3317# VGND 1.92f $ **FLOATING
C218 a_12056_3689# VGND 0.736f $ **FLOATING
C219 a_12231_3615# VGND 1.54f $ **FLOATING
C220 a_11491_3689# VGND 0.714f $ **FLOATING
C221 a_11709_3285# VGND 0.653f $ **FLOATING
C222 a_11141_3317# VGND 1.57f $ **FLOATING
C223 a_10975_3317# VGND 1.92f $ **FLOATING
C224 a_10523_3427# VGND 0.485f $ **FLOATING
C225 a_10331_3671# VGND 0.478f $ **FLOATING
C226 a_9414_3311# VGND 0.259f $ **FLOATING
C227 a_10011_3530# VGND 0.524f $ **FLOATING
C228 _027_ VGND 1.02f $ **FLOATING
C229 a_8782_3311# VGND 0.653f $ **FLOATING
C230 a_8851_3285# VGND 0.714f $ **FLOATING
C231 a_8656_3427# VGND 1.57f $ **FLOATING
C232 a_8695_3553# VGND 1.92f $ **FLOATING
C233 a_8378_3443# VGND 0.736f $ **FLOATING
C234 a_8175_3285# VGND 0.971f $ **FLOATING
C235 a_6791_3530# VGND 0.524f $ **FLOATING
C236 a_3519_3311# VGND 0.553f $ **FLOATING
C237 a_3413_3311# VGND 0.794f $ **FLOATING
C238 a_3177_3311# VGND 0.788f $ **FLOATING
C239 a_15741_3855# VGND 0.824f $ **FLOATING
C240 a_14085_3855# VGND 0.824f $ **FLOATING
C241 a_11808_3855# VGND 0.824f $ **FLOATING
C242 a_10313_3855# VGND 0.824f $ **FLOATING
C243 a_15763_4117# VGND 1.18f $ **FLOATING
C244 a_14107_4117# VGND 1.18f $ **FLOATING
C245 a_11812_4105# VGND 1.18f $ **FLOATING
C246 a_10335_4117# VGND 1.18f $ **FLOATING
C247 a_8877_3829# VGND 0.607f $ **FLOATING
C248 _222_ VGND 1.47f $ **FLOATING
C249 a_6907_4221# VGND 0.168f $ **FLOATING
C250 a_6704_3855# VGND 0.259f $ **FLOATING
C251 a_18755_3829# VGND 0.698f $ **FLOATING
C252 a_18293_4020# VGND 0.524f $ **FLOATING
C253 a_17332_3829# VGND 1.98f $ **FLOATING
C254 a_15575_3855# VGND 1.46f $ **FLOATING
C255 a_13919_3855# VGND 1.46f $ **FLOATING
C256 a_12547_4007# VGND 1.46f $ **FLOATING
C257 net71 VGND 9.75f $ **FLOATING
C258 a_10147_3855# VGND 1.46f $ **FLOATING
C259 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd VGND 14.4f $ **FLOATING
C260 a_9287_3829# VGND 1.2f $ **FLOATING
C261 a_8448_4007# VGND 0.59f $ **FLOATING
C262 a_7364_3855# VGND 0.736f $ **FLOATING
C263 a_7539_3829# VGND 0.971f $ **FLOATING
C264 a_6799_3855# VGND 0.714f $ **FLOATING
C265 a_7017_4097# VGND 0.653f $ **FLOATING
C266 a_6449_3855# VGND 1.57f $ **FLOATING
C267 _046_ VGND 1.12f $ **FLOATING
C268 a_6283_3855# VGND 1.92f $ **FLOATING
C269 a_3601_3855# VGND 0.23f $ **FLOATING
C270 a_4111_4221# VGND 0.609f $ **FLOATING
C271 a_4279_4123# VGND 0.817f $ **FLOATING
C272 a_3686_4221# VGND 0.626f $ **FLOATING
C273 a_3854_3967# VGND 0.581f $ **FLOATING
C274 a_3413_3855# VGND 1.43f $ **FLOATING
C275 net56 VGND 1.06f $ **FLOATING
C276 a_3247_3855# VGND 1.81f $ **FLOATING
C277 net52 VGND 0.786f $ **FLOATING
C278 res1_n VGND 1.1f $ **FLOATING
C279 a_1761_3855# VGND 0.23f $ **FLOATING
C280 a_2271_4221# VGND 0.609f $ **FLOATING
C281 a_2439_4123# VGND 0.817f $ **FLOATING
C282 a_1846_4221# VGND 0.626f $ **FLOATING
C283 a_2014_3967# VGND 0.581f $ **FLOATING
C284 a_1573_3855# VGND 1.43f $ **FLOATING
C285 a_1407_3855# VGND 1.81f $ **FLOATING
C286 net53 VGND 0.747f $ **FLOATING
C287 a_17695_4399# VGND 1.18f $ **FLOATING
C288 a_16129_4399# VGND 0.253f $ **FLOATING
C289 a_14296_4399# VGND 1.18f $ **FLOATING
C290 a_17673_4719# VGND 0.824f $ **FLOATING
C291 a_17507_4399# VGND 1.46f $ **FLOATING
C292 a_16863_4719# VGND 0.275f $ **FLOATING
C293 _006_ VGND 2.68f $ **FLOATING
C294 a_15031_4373# VGND 1.46f $ **FLOATING
C295 a_14292_4719# VGND 0.824f $ **FLOATING
C296 a_12427_4399# VGND 0.168f $ **FLOATING
C297 a_11255_4399# VGND 0.19f $ **FLOATING
C298 a_12224_4765# VGND 0.259f $ **FLOATING
C299 a_9765_4399# VGND 0.23f $ **FLOATING
C300 _202_ VGND 1.7f $ **FLOATING
C301 _145_ VGND 4.98f $ **FLOATING
C302 a_6631_4399# VGND 0.168f $ **FLOATING
C303 a_6428_4765# VGND 0.259f $ **FLOATING
C304 a_4515_4399# VGND 0.168f $ **FLOATING
C305 a_4312_4765# VGND 0.259f $ **FLOATING
C306 net1 VGND 1.26f $ **FLOATING
C307 a_17017_4399# VGND 0.597f $ **FLOATING
C308 a_16298_4719# VGND 0.55f $ **FLOATING
C309 net65 VGND 1.29f $ **FLOATING
C310 a_12884_4777# VGND 0.736f $ **FLOATING
C311 a_13059_4703# VGND 1.54f $ **FLOATING
C312 a_12319_4777# VGND 0.714f $ **FLOATING
C313 a_12537_4373# VGND 0.653f $ **FLOATING
C314 a_11969_4405# VGND 1.57f $ **FLOATING
C315 _005_ VGND 1.26f $ **FLOATING
C316 a_11803_4405# VGND 1.92f $ **FLOATING
C317 a_11478_4373# VGND 0.552f $ **FLOATING
C318 a_11119_4373# VGND 0.629f $ **FLOATING
C319 a_10275_4399# VGND 0.609f $ **FLOATING
C320 a_10443_4373# VGND 0.817f $ **FLOATING
C321 a_9850_4399# VGND 0.626f $ **FLOATING
C322 a_10018_4373# VGND 0.581f $ **FLOATING
C323 a_9577_4405# VGND 1.43f $ **FLOATING
C324 net57 VGND 2.6f $ **FLOATING
C325 a_9411_4405# VGND 1.81f $ **FLOATING
C326 net55 VGND 2.3f $ **FLOATING
C327 a_8879_4438# VGND 0.59f $ **FLOATING
C328 a_8625_4438# VGND 0.607f $ **FLOATING
C329 a_8155_4737# VGND 0.56f $ **FLOATING
C330 a_7088_4777# VGND 0.736f $ **FLOATING
C331 a_7263_4703# VGND 0.971f $ **FLOATING
C332 a_6523_4777# VGND 0.714f $ **FLOATING
C333 a_6741_4373# VGND 0.653f $ **FLOATING
C334 a_6173_4405# VGND 1.57f $ **FLOATING
C335 a_6007_4405# VGND 1.92f $ **FLOATING
C336 a_4972_4777# VGND 0.736f $ **FLOATING
C337 a_5147_4703# VGND 0.971f $ **FLOATING
C338 a_4407_4777# VGND 0.714f $ **FLOATING
C339 a_4625_4373# VGND 0.653f $ **FLOATING
C340 a_4057_4405# VGND 1.57f $ **FLOATING
C341 a_3891_4405# VGND 1.92f $ **FLOATING
C342 a_855_4399# VGND 0.524f $ **FLOATING
C343 a_17121_4943# VGND 0.824f $ **FLOATING
C344 a_16311_4943# VGND 0.275f $ **FLOATING
C345 a_14453_4943# VGND 0.824f $ **FLOATING
C346 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref VGND 8.79f $ **FLOATING
C347 a_18719_5193# VGND 0.388f $ **FLOATING
C348 a_17143_5205# VGND 1.18f $ **FLOATING
C349 a_16955_4943# VGND 1.46f $ **FLOATING
C350 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref VGND 2.27f $ **FLOATING
C351 a_16465_5193# VGND 0.597f $ **FLOATING
C352 a_15943_4943# VGND 0.648f $ **FLOATING
C353 a_11808_4943# VGND 0.824f $ **FLOATING
C354 a_10883_4943# VGND 0.171f $ **FLOATING
C355 a_14475_5205# VGND 1.18f $ **FLOATING
C356 a_11812_5193# VGND 1.18f $ **FLOATING
C357 _004_ VGND 1.51f $ **FLOATING
C358 a_9391_5309# VGND 0.168f $ **FLOATING
C359 a_9188_4943# VGND 0.259f $ **FLOATING
C360 a_14287_4943# VGND 1.46f $ **FLOATING
C361 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd VGND 5.24f $ **FLOATING
C362 a_13611_4917# VGND 1.2f $ **FLOATING
C363 a_12547_5095# VGND 1.46f $ **FLOATING
C364 a_11056_5193# VGND 0.546f $ **FLOATING
C365 _156_ VGND 2.01f $ **FLOATING
C366 _155_ VGND 1.47f $ **FLOATING
C367 a_9848_4943# VGND 0.736f $ **FLOATING
C368 a_10023_4917# VGND 0.971f $ **FLOATING
C369 a_9283_4943# VGND 0.714f $ **FLOATING
C370 a_9501_5185# VGND 0.653f $ **FLOATING
C371 a_8933_4943# VGND 1.57f $ **FLOATING
C372 a_8767_4943# VGND 1.92f $ **FLOATING
C373 a_7313_4917# VGND 0.607f $ **FLOATING
C374 _045_ VGND 1.13f $ **FLOATING
C375 a_4055_5309# VGND 0.168f $ **FLOATING
C376 a_3852_4943# VGND 0.259f $ **FLOATING
C377 a_7815_4917# VGND 1.2f $ **FLOATING
C378 a_6884_5095# VGND 0.59f $ **FLOATING
C379 _221_ VGND 0.73f $ **FLOATING
C380 a_6515_5108# VGND 0.524f $ **FLOATING
C381 a_5423_4917# VGND 1.2f $ **FLOATING
C382 a_4512_4943# VGND 0.736f $ **FLOATING
C383 a_4687_4917# VGND 0.971f $ **FLOATING
C384 a_3947_4943# VGND 0.714f $ **FLOATING
C385 a_4165_5185# VGND 0.653f $ **FLOATING
C386 a_3597_4943# VGND 1.57f $ **FLOATING
C387 a_3431_4943# VGND 1.92f $ **FLOATING
C388 a_16315_5487# VGND 1.18f $ **FLOATING
C389 a_15591_5487# VGND 0.388f $ **FLOATING
C390 a_13928_5487# VGND 1.18f $ **FLOATING
C391 a_16293_5807# VGND 0.824f $ **FLOATING
C392 a_16127_5487# VGND 1.46f $ **FLOATING
C393 a_14663_5461# VGND 1.46f $ **FLOATING
C394 a_13924_5807# VGND 0.824f $ **FLOATING
C395 a_13463_5807# VGND 0.275f $ **FLOATING
C396 a_17783_5487# VGND 2.1f $ **FLOATING
C397 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd VGND 6.51f $ **FLOATING
C398 a_13326_5719# VGND 0.597f $ **FLOATING
C399 a_12447_5540# VGND 0.732f $ **FLOATING
C400 net15 VGND 19.2f $ **FLOATING
C401 _147_ VGND 2.69f $ **FLOATING
C402 _146_ VGND 4.76f $ **FLOATING
C403 _153_ VGND 4.25f $ **FLOATING
C404 _007_ VGND 1.4f $ **FLOATING
C405 a_8287_5487# VGND 0.168f $ **FLOATING
C406 a_8084_5853# VGND 0.259f $ **FLOATING
C407 a_5085_5487# VGND 0.203f $ **FLOATING
C408 _026_ VGND 1.58f $ **FLOATING
C409 a_4588_5807# VGND 0.205f $ **FLOATING
C410 _025_ VGND 1.21f $ **FLOATING
C411 a_2859_5487# VGND 0.168f $ **FLOATING
C412 a_2656_5853# VGND 0.259f $ **FLOATING
C413 a_12596_5461# VGND 0.719f $ **FLOATING
C414 a_11975_5461# VGND 0.988f $ **FLOATING
C415 a_11467_5825# VGND 0.56f $ **FLOATING
C416 a_11053_5719# VGND 0.502f $ **FLOATING
C417 a_10441_5785# VGND 0.607f $ **FLOATING
C418 a_10012_5719# VGND 0.59f $ **FLOATING
C419 _157_ VGND 0.878f $ **FLOATING
C420 a_8744_5865# VGND 0.736f $ **FLOATING
C421 a_8919_5791# VGND 0.971f $ **FLOATING
C422 a_8179_5865# VGND 0.714f $ **FLOATING
C423 a_8397_5461# VGND 0.653f $ **FLOATING
C424 a_7829_5493# VGND 1.57f $ **FLOATING
C425 a_7663_5493# VGND 1.92f $ **FLOATING
C426 a_6559_5487# VGND 1.2f $ **FLOATING
C427 a_6247_5461# VGND 0.788f $ **FLOATING
C428 a_5989_5461# VGND 0.794f $ **FLOATING
C429 a_5893_5719# VGND 0.553f $ **FLOATING
C430 a_4956_5461# VGND 0.655f $ **FLOATING
C431 net59 VGND 1.35f $ **FLOATING
C432 a_4362_5603# VGND 0.443f $ **FLOATING
C433 a_4219_5461# VGND 0.65f $ **FLOATING
C434 a_3316_5865# VGND 0.736f $ **FLOATING
C435 a_3491_5791# VGND 1.13f $ **FLOATING
C436 a_2751_5865# VGND 0.714f $ **FLOATING
C437 a_2969_5461# VGND 0.653f $ **FLOATING
C438 a_2401_5493# VGND 1.57f $ **FLOATING
C439 a_2235_5493# VGND 1.92f $ **FLOATING
C440 _142_ VGND 1.59f $ **FLOATING
C441 a_17599_6031# VGND 0.424f $ **FLOATING
C442 a_16109_6031# VGND 0.824f $ **FLOATING
C443 a_14453_6031# VGND 0.824f $ **FLOATING
C444 a_13551_6031# VGND 0.186f $ **FLOATING
C445 a_17862_6281# VGND 0.171f $ **FLOATING
C446 a_16131_6293# VGND 1.18f $ **FLOATING
C447 a_14475_6293# VGND 1.18f $ **FLOATING
C448 a_12997_6031# VGND 0.277f $ **FLOATING
C449 _063_ VGND 2.34f $ **FLOATING
C450 a_13769_6296# VGND 0.538f $ **FLOATING
C451 a_10403_6397# VGND 0.168f $ **FLOATING
C452 a_10200_6031# VGND 0.259f $ **FLOATING
C453 a_9245_6005# VGND 0.607f $ **FLOATING
C454 a_18735_6059# VGND 0.56f $ **FLOATING
C455 a_15943_6031# VGND 1.46f $ **FLOATING
C456 a_14287_6031# VGND 1.46f $ **FLOATING
C457 a_13705_6353# VGND 0.645f $ **FLOATING
C458 net5 VGND 4.35f $ **FLOATING
C459 a_12777_6005# VGND 0.758f $ **FLOATING
C460 a_12275_6281# VGND 0.642f $ **FLOATING
C461 a_11679_6183# VGND 0.56f $ **FLOATING
C462 a_10860_6031# VGND 0.736f $ **FLOATING
C463 a_11035_6005# VGND 0.971f $ **FLOATING
C464 a_10295_6031# VGND 0.714f $ **FLOATING
C465 a_10513_6273# VGND 0.653f $ **FLOATING
C466 a_9945_6031# VGND 1.57f $ **FLOATING
C467 a_9779_6031# VGND 1.92f $ **FLOATING
C468 _028_ VGND 1.3f $ **FLOATING
C469 a_7313_6005# VGND 0.607f $ **FLOATING
C470 a_5361_6281# VGND 0.203f $ **FLOATING
C471 _199_ VGND 1.35f $ **FLOATING
C472 _201_ VGND 1.67f $ **FLOATING
C473 a_4617_6281# VGND 0.212f $ **FLOATING
C474 _198_ VGND 1.34f $ **FLOATING
C475 a_8816_6183# VGND 0.59f $ **FLOATING
C476 _203_ VGND 0.73f $ **FLOATING
C477 a_8447_6196# VGND 0.524f $ **FLOATING
C478 a_6884_6183# VGND 0.59f $ **FLOATING
C479 _220_ VGND 0.73f $ **FLOATING
C480 a_6515_6196# VGND 0.524f $ **FLOATING
C481 _136_ VGND 3.01f $ **FLOATING
C482 a_6059_6005# VGND 0.698f $ **FLOATING
C483 a_5232_6005# VGND 0.655f $ **FLOATING
C484 _200_ VGND 2.21f $ **FLOATING
C485 a_4075_6031# VGND 0.619f $ **FLOATING
C486 a_17695_6575# VGND 1.18f $ **FLOATING
C487 a_16609_6575# VGND 0.336f $ **FLOATING
C488 a_14567_6575# VGND 1.18f $ **FLOATING
C489 a_17673_6895# VGND 0.824f $ **FLOATING
C490 a_17507_6575# VGND 1.46f $ **FLOATING
C491 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd VGND 11.7f $ **FLOATING
C492 a_16170_6895# VGND 0.54f $ **FLOATING
C493 a_14545_6895# VGND 0.824f $ **FLOATING
C494 a_14379_6575# VGND 1.46f $ **FLOATING
C495 a_12591_6895# VGND 0.509f $ **FLOATING
C496 a_10141_6575# VGND 0.238f $ **FLOATING
C497 a_6631_6575# VGND 0.168f $ **FLOATING
C498 a_6428_6941# VGND 0.259f $ **FLOATING
C499 _024_ VGND 1.49f $ **FLOATING
C500 a_1769_6895# VGND 0.171f $ **FLOATING
C501 net68 VGND 10.6f $ **FLOATING
C502 net4 VGND 6.1f $ **FLOATING
C503 a_13963_6896# VGND 0.641f $ **FLOATING
C504 a_13599_6807# VGND 0.673f $ **FLOATING
C505 a_12047_6835# VGND 1.2f $ **FLOATING
C506 _062_ VGND 7.35f $ **FLOATING
C507 a_11339_6575# VGND 0.508f $ **FLOATING
C508 a_11159_6575# VGND 0.604f $ **FLOATING
C509 _112_ VGND 6.88f $ **FLOATING
C510 a_8022_6575# VGND 4.03f $ **FLOATING
C511 a_7088_6953# VGND 0.736f $ **FLOATING
C512 a_7263_6879# VGND 0.971f $ **FLOATING
C513 a_6523_6953# VGND 0.714f $ **FLOATING
C514 a_6741_6549# VGND 0.653f $ **FLOATING
C515 a_6173_6581# VGND 1.57f $ **FLOATING
C516 _044_ VGND 1.15f $ **FLOATING
C517 a_6007_6581# VGND 1.92f $ **FLOATING
C518 clknet_2_1__leaf_clk VGND 15.6f $ **FLOATING
C519 _196_ VGND 0.876f $ **FLOATING
C520 a_3479_6807# VGND 0.619f $ **FLOATING
C521 _197_ VGND 0.722f $ **FLOATING
C522 a_3111_6794# VGND 0.524f $ **FLOATING
C523 a_2751_6549# VGND 0.788f $ **FLOATING
C524 a_2493_6549# VGND 0.794f $ **FLOATING
C525 a_2397_6807# VGND 0.553f $ **FLOATING
C526 net61 VGND 0.732f $ **FLOATING
C527 a_1551_6807# VGND 0.546f $ **FLOATING
C528 a_17121_7119# VGND 0.824f $ **FLOATING
C529 a_15304_7119# VGND 0.824f $ **FLOATING
C530 a_17143_7381# VGND 1.18f $ **FLOATING
C531 a_12851_7119# VGND 0.398f $ **FLOATING
C532 a_12493_7119# VGND 0.155f $ **FLOATING
C533 a_15308_7369# VGND 1.18f $ **FLOATING
C534 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref VGND 16.1f $ **FLOATING
C535 a_13845_7369# VGND 1.19f $ **FLOATING
C536 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd VGND 4.26f $ **FLOATING
C537 a_13101_7369# VGND 0.171f $ **FLOATING
C538 a_11437_7369# VGND 0.253f $ **FLOATING
C539 _008_ VGND 1.73f $ **FLOATING
C540 a_8481_7369# VGND 0.206f $ **FLOATING
C541 a_7221_7093# VGND 0.607f $ **FLOATING
C542 a_4071_7369# VGND 0.253f $ **FLOATING
C543 _195_ VGND 1.01f $ **FLOATING
C544 a_1479_7485# VGND 0.168f $ **FLOATING
C545 a_1276_7119# VGND 0.259f $ **FLOATING
C546 a_18763_7271# VGND 0.56f $ **FLOATING
C547 a_16955_7119# VGND 1.46f $ **FLOATING
C548 net67 VGND 22.4f $ **FLOATING
C549 a_16043_7271# VGND 1.46f $ **FLOATING
C550 net14 VGND 26.9f $ **FLOATING
C551 _144_ VGND 6.39f $ **FLOATING
C552 a_13551_7119# VGND 0.524f $ **FLOATING
C553 _111_ VGND 3.62f $ **FLOATING
C554 a_12493_7369# VGND 0.822f $ **FLOATING
C555 _110_ VGND 2.83f $ **FLOATING
C556 a_12127_7093# VGND 1.43f $ **FLOATING
C557 a_11606_7119# VGND 0.55f $ **FLOATING
C558 a_10625_7352# VGND 0.696f $ **FLOATING
C559 a_10147_7119# VGND 0.788f $ **FLOATING
C560 a_10294_7093# VGND 0.795f $ **FLOATING
C561 _158_ VGND 1.23f $ **FLOATING
C562 a_8399_7369# VGND 0.804f $ **FLOATING
C563 ts.ts_ctrl.temp_ctr\[18\] VGND 6.16f $ **FLOATING
C564 a_6792_7271# VGND 0.59f $ **FLOATING
C565 a_4986_7119# VGND 4.03f $ **FLOATING
C566 a_3853_7093# VGND 0.55f $ **FLOATING
C567 a_1936_7119# VGND 0.736f $ **FLOATING
C568 a_2111_7093# VGND 1.13f $ **FLOATING
C569 a_1371_7119# VGND 0.714f $ **FLOATING
C570 a_1589_7361# VGND 0.653f $ **FLOATING
C571 a_1021_7119# VGND 1.57f $ **FLOATING
C572 _009_ VGND 1.28f $ **FLOATING
C573 a_855_7119# VGND 1.92f $ **FLOATING
C574 a_18691_7663# VGND 0.381f $ **FLOATING
C575 a_18243_7663# VGND 0.381f $ **FLOATING
C576 a_16775_7663# VGND 1.18f $ **FLOATING
C577 a_18243_7983# VGND 0.554f $ **FLOATING
C578 a_16753_7983# VGND 0.824f $ **FLOATING
C579 a_15321_7663# VGND 0.336f $ **FLOATING
C580 a_13183_7663# VGND 1.23f $ **FLOATING
C581 a_12691_7663# VGND 0.203f $ **FLOATING
C582 a_12181_7663# VGND 0.171f $ **FLOATING
C583 a_8573_7663# VGND 0.206f $ **FLOATING
C584 a_7929_7663# VGND 0.206f $ **FLOATING
C585 a_16587_7663# VGND 1.46f $ **FLOATING
C586 _060_ VGND 2.94f $ **FLOATING
C587 a_14882_7983# VGND 0.54f $ **FLOATING
C588 a_13601_7983# VGND 0.309f $ **FLOATING
C589 a_13183_7983# VGND 0.43f $ **FLOATING
C590 a_11931_7983# VGND 0.398f $ **FLOATING
C591 a_11573_7983# VGND 0.155f $ **FLOATING
C592 a_6447_7663# VGND 0.168f $ **FLOATING
C593 a_1769_7663# VGND 0.238f $ **FLOATING
C594 a_6244_8029# VGND 0.259f $ **FLOATING
C595 _160_ VGND 0.997f $ **FLOATING
C596 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd VGND 7.55f $ **FLOATING
C597 a_16187_7895# VGND 0.56f $ **FLOATING
C598 net6 VGND 5.27f $ **FLOATING
C599 a_12597_7663# VGND 0.655f $ **FLOATING
C600 _113_ VGND 3.94f $ **FLOATING
C601 _096_ VGND 3.74f $ **FLOATING
C602 a_11573_7663# VGND 0.822f $ **FLOATING
C603 _058_ VGND 6.52f $ **FLOATING
C604 a_11207_7637# VGND 1.43f $ **FLOATING
C605 a_8491_7663# VGND 0.804f $ **FLOATING
C606 ts.ts_ctrl.temp_ctr\[17\] VGND 7.13f $ **FLOATING
C607 a_7847_7663# VGND 0.804f $ **FLOATING
C608 ts.ts_ctrl.temp_ctr\[19\] VGND 5.02f $ **FLOATING
C609 a_6904_8041# VGND 0.736f $ **FLOATING
C610 a_7079_7967# VGND 0.971f $ **FLOATING
C611 a_6339_8041# VGND 0.714f $ **FLOATING
C612 a_6557_7637# VGND 0.653f $ **FLOATING
C613 a_5989_7669# VGND 1.57f $ **FLOATING
C614 _029_ VGND 1.06f $ **FLOATING
C615 a_5823_7669# VGND 1.92f $ **FLOATING
C616 a_5455_7663# VGND 0.524f $ **FLOATING
C617 _204_ VGND 1.44f $ **FLOATING
C618 a_17121_8207# VGND 0.824f $ **FLOATING
C619 a_15304_8207# VGND 0.824f $ **FLOATING
C620 a_14471_8207# VGND 0.509f $ **FLOATING
C621 a_14024_8207# VGND 0.238f $ **FLOATING
C622 a_13834_8207# VGND 0.217f $ **FLOATING
C623 _150_ VGND 3.55f $ **FLOATING
C624 _151_ VGND 3.41f $ **FLOATING
C625 a_17143_8469# VGND 1.18f $ **FLOATING
C626 a_15308_8457# VGND 1.18f $ **FLOATING
C627 a_12631_8457# VGND 0.388f $ **FLOATING
C628 _125_ VGND 1.41f $ **FLOATING
C629 _115_ VGND 2.29f $ **FLOATING
C630 _124_ VGND 0.627f $ **FLOATING
C631 a_11610_8457# VGND 0.191f $ **FLOATING
C632 ts.o_res\[17\] VGND 3.75f $ **FLOATING
C633 a_8809_8534# VGND 0.607f $ **FLOATING
C634 ts.o_res\[18\] VGND 4.19f $ **FLOATING
C635 a_7521_8534# VGND 0.607f $ **FLOATING
C636 a_6209_8181# VGND 0.607f $ **FLOATING
C637 a_3871_8573# VGND 0.168f $ **FLOATING
C638 a_3668_8207# VGND 0.259f $ **FLOATING
C639 a_18763_8359# VGND 0.56f $ **FLOATING
C640 a_16955_8207# VGND 1.46f $ **FLOATING
C641 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd VGND 4.27f $ **FLOATING
C642 a_16043_8359# VGND 1.46f $ **FLOATING
C643 a_13643_8207# VGND 0.893f $ **FLOATING
C644 net7 VGND 6.5f $ **FLOATING
C645 a_13183_8207# VGND 0.524f $ **FLOATING
C646 _149_ VGND 3.65f $ **FLOATING
C647 a_12079_8457# VGND 0.702f $ **FLOATING
C648 a_11435_8207# VGND 0.847f $ **FLOATING
C649 _122_ VGND 3.74f $ **FLOATING
C650 _123_ VGND 2.04f $ **FLOATING
C651 a_9063_8534# VGND 0.59f $ **FLOATING
C652 a_7775_8534# VGND 0.59f $ **FLOATING
C653 a_5780_8359# VGND 0.59f $ **FLOATING
C654 a_4328_8207# VGND 0.736f $ **FLOATING
C655 a_4503_8181# VGND 0.971f $ **FLOATING
C656 a_3763_8207# VGND 0.714f $ **FLOATING
C657 a_3981_8449# VGND 0.653f $ **FLOATING
C658 a_3413_8207# VGND 1.57f $ **FLOATING
C659 a_3247_8207# VGND 1.92f $ **FLOATING
C660 a_1775_8457# VGND 0.238f $ **FLOATING
C661 _161_ VGND 0.807f $ **FLOATING
C662 a_17695_8751# VGND 1.18f $ **FLOATING
C663 a_16793_8751# VGND 0.336f $ **FLOATING
C664 a_14852_8751# VGND 0.14f $ **FLOATING
C665 a_14500_8751# VGND 0.171f $ **FLOATING
C666 a_17673_9071# VGND 0.824f $ **FLOATING
C667 a_17507_8751# VGND 1.46f $ **FLOATING
C668 a_16354_9071# VGND 0.54f $ **FLOATING
C669 a_14418_9071# VGND 0.482f $ **FLOATING
C670 a_9687_8751# VGND 0.333f $ **FLOATING
C671 a_6447_8751# VGND 0.168f $ **FLOATING
C672 a_4713_8751# VGND 0.238f $ **FLOATING
C673 a_6244_9117# VGND 0.259f $ **FLOATING
C674 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd VGND 6.64f $ **FLOATING
C675 a_14584_8751# VGND 1.37f $ **FLOATING
C676 _064_ VGND 2.29f $ **FLOATING
C677 a_13731_8751# VGND 0.508f $ **FLOATING
C678 a_13551_8751# VGND 0.604f $ **FLOATING
C679 a_11435_8864# VGND 0.619f $ **FLOATING
C680 ts.ts_ctrl.state\[1\] VGND 11.5f $ **FLOATING
C681 a_10975_8864# VGND 0.619f $ **FLOATING
C682 a_9770_8751# VGND 0.723f $ **FLOATING
C683 ts.ts_ctrl.state\[0\] VGND 13.5f $ **FLOATING
C684 a_8235_8790# VGND 0.59f $ **FLOATING
C685 ts.o_res\[19\] VGND 4.17f $ **FLOATING
C686 a_7981_8790# VGND 0.607f $ **FLOATING
C687 a_6904_9129# VGND 0.736f $ **FLOATING
C688 a_7079_9055# VGND 0.971f $ **FLOATING
C689 a_6339_9129# VGND 0.714f $ **FLOATING
C690 a_6557_8725# VGND 0.653f $ **FLOATING
C691 a_5989_8757# VGND 1.57f $ **FLOATING
C692 _030_ VGND 1.1f $ **FLOATING
C693 a_5823_8757# VGND 1.92f $ **FLOATING
C694 a_5363_8751# VGND 0.524f $ **FLOATING
C695 _205_ VGND 1.01f $ **FLOATING
C696 _023_ VGND 1.32f $ **FLOATING
C697 ts.ts_ctrl.temp_ctr\[2\] VGND 8.98f $ **FLOATING
C698 a_1479_8751# VGND 0.168f $ **FLOATING
C699 a_1276_9117# VGND 0.259f $ **FLOATING
C700 a_4126_8983# VGND 0.759f $ **FLOATING
C701 _194_ VGND 4.79f $ **FLOATING
C702 _193_ VGND 1f $ **FLOATING
C703 a_2755_8983# VGND 0.56f $ **FLOATING
C704 a_1936_9129# VGND 0.736f $ **FLOATING
C705 a_2111_9055# VGND 0.971f $ **FLOATING
C706 a_1371_9129# VGND 0.714f $ **FLOATING
C707 net16 VGND 18.8f $ **FLOATING
C708 a_1589_8725# VGND 0.653f $ **FLOATING
C709 a_1021_8757# VGND 1.57f $ **FLOATING
C710 _010_ VGND 1.48f $ **FLOATING
C711 a_855_8757# VGND 1.92f $ **FLOATING
C712 clknet_2_0__leaf_clk VGND 15.5f $ **FLOATING
C713 a_17599_9295# VGND 0.275f $ **FLOATING
C714 a_15948_9295# VGND 0.824f $ **FLOATING
C715 a_14195_9295# VGND 0.594f $ **FLOATING
C716 _139_ VGND 10.4f $ **FLOATING
C717 _148_ VGND 2.75f $ **FLOATING
C718 a_15952_9545# VGND 1.18f $ **FLOATING
C719 a_14907_9545# VGND 0.399f $ **FLOATING
C720 a_14445_9545# VGND 0.384f $ **FLOATING
C721 a_14195_9545# VGND 0.388f $ **FLOATING
C722 _108_ VGND 1.8f $ **FLOATING
C723 _105_ VGND 0.745f $ **FLOATING
C724 a_11877_9545# VGND 0.214f $ **FLOATING
C725 a_11793_9545# VGND 0.167f $ **FLOATING
C726 a_11150_9545# VGND 0.191f $ **FLOATING
C727 _107_ VGND 1.28f $ **FLOATING
C728 a_10405_9545# VGND 0.214f $ **FLOATING
C729 a_10321_9545# VGND 0.167f $ **FLOATING
C730 a_9669_9545# VGND 0.214f $ **FLOATING
C731 a_9585_9545# VGND 0.167f $ **FLOATING
C732 a_8877_9269# VGND 0.607f $ **FLOATING
C733 ts.ts_ctrl.temp_ctr\[16\] VGND 4.59f $ **FLOATING
C734 a_6631_9661# VGND 0.168f $ **FLOATING
C735 a_6428_9295# VGND 0.259f $ **FLOATING
C736 a_18763_9447# VGND 0.56f $ **FLOATING
C737 _143_ VGND 9.19f $ **FLOATING
C738 _141_ VGND 3.77f $ **FLOATING
C739 a_17753_9545# VGND 0.597f $ **FLOATING
C740 _140_ VGND 9f $ **FLOATING
C741 _098_ VGND 8.99f $ **FLOATING
C742 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref VGND 5f $ **FLOATING
C743 a_16687_9447# VGND 1.46f $ **FLOATING
C744 a_14717_9545# VGND 1.44f $ **FLOATING
C745 _134_ VGND 1.51f $ **FLOATING
C746 a_12449_9301# VGND 0.665f $ **FLOATING
C747 a_11711_9295# VGND 0.972f $ **FLOATING
C748 ts.ts_ctrl.temp_ctr\[1\] VGND 5.03f $ **FLOATING
C749 _104_ VGND 0.811f $ **FLOATING
C750 a_10975_9295# VGND 0.847f $ **FLOATING
C751 _109_ VGND 2.19f $ **FLOATING
C752 a_10239_9295# VGND 0.972f $ **FLOATING
C753 ts.o_res\[1\] VGND 3.95f $ **FLOATING
C754 _106_ VGND 1.69f $ **FLOATING
C755 a_9503_9295# VGND 0.972f $ **FLOATING
C756 ts.ts_ctrl.temp_ctr\[0\] VGND 6.19f $ **FLOATING
C757 _091_ VGND 1.12f $ **FLOATING
C758 a_8448_9447# VGND 0.59f $ **FLOATING
C759 a_7088_9295# VGND 0.736f $ **FLOATING
C760 a_7263_9269# VGND 0.971f $ **FLOATING
C761 a_6523_9295# VGND 0.714f $ **FLOATING
C762 net17 VGND 20f $ **FLOATING
C763 a_6741_9537# VGND 0.653f $ **FLOATING
C764 a_6173_9295# VGND 1.57f $ **FLOATING
C765 a_6007_9295# VGND 1.92f $ **FLOATING
C766 _163_ VGND 0.894f $ **FLOATING
C767 a_3299_9269# VGND 0.698f $ **FLOATING
C768 a_2451_9323# VGND 0.56f $ **FLOATING
C769 a_17603_9839# VGND 1.18f $ **FLOATING
C770 a_17034_9839# VGND 0.171f $ **FLOATING
C771 a_17581_10159# VGND 0.824f $ **FLOATING
C772 a_17415_9839# VGND 1.46f $ **FLOATING
C773 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd VGND 6.89f $ **FLOATING
C774 a_16771_10159# VGND 0.424f $ **FLOATING
C775 _100_ VGND 2.32f $ **FLOATING
C776 a_16127_10159# VGND 0.277f $ **FLOATING
C777 _097_ VGND 2.4f $ **FLOATING
C778 _061_ VGND 11.9f $ **FLOATING
C779 _065_ VGND 9.68f $ **FLOATING
C780 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd VGND 6.71f $ **FLOATING
C781 _099_ VGND 3.95f $ **FLOATING
C782 _095_ VGND 5.34f $ **FLOATING
C783 a_14937_9955# VGND 0.828f $ **FLOATING
C784 a_14986_9849# VGND 0.812f $ **FLOATING
C785 _135_ VGND 1.01f $ **FLOATING
C786 _089_ VGND 3.21f $ **FLOATING
C787 a_14177_9839# VGND 0.673f $ **FLOATING
C788 ts.ts_core.i_precharge_n VGND 4.5f $ **FLOATING
C789 a_14011_9839# VGND 0.641f $ **FLOATING
C790 a_13503_10145# VGND 0.604f $ **FLOATING
C791 a_13327_9813# VGND 0.508f $ **FLOATING
C792 a_12952_10071# VGND 0.488f $ **FLOATING
C793 a_10229_9839# VGND 0.206f $ **FLOATING
C794 a_9045_9839# VGND 0.253f $ **FLOATING
C795 _093_ VGND 2.22f $ **FLOATING
C796 a_12679_10071# VGND 0.601f $ **FLOATING
C797 a_12157_9813# VGND 0.713f $ **FLOATING
C798 a_10977_9955# VGND 0.665f $ **FLOATING
C799 _092_ VGND 1.24f $ **FLOATING
C800 _126_ VGND 1.48f $ **FLOATING
C801 _133_ VGND 2.95f $ **FLOATING
C802 a_10147_9839# VGND 0.804f $ **FLOATING
C803 ts.o_res\[3\] VGND 4.42f $ **FLOATING
C804 a_9597_9955# VGND 0.665f $ **FLOATING
C805 _128_ VGND 1.65f $ **FLOATING
C806 _130_ VGND 0.709f $ **FLOATING
C807 _043_ VGND 1.16f $ **FLOATING
C808 a_9214_10159# VGND 0.55f $ **FLOATING
C809 ts.ts_ctrl.temp_ctr\[3\] VGND 6.61f $ **FLOATING
C810 _087_ VGND 5.87f $ **FLOATING
C811 a_7286_9839# VGND 4.03f $ **FLOATING
C812 _219_ VGND 1.6f $ **FLOATING
C813 a_6515_10058# VGND 0.524f $ **FLOATING
C814 a_3431_9839# VGND 0.698f $ **FLOATING
C815 _171_ VGND 0.663f $ **FLOATING
C816 a_2787_10205# VGND 0.729f $ **FLOATING
C817 _162_ VGND 2.08f $ **FLOATING
C818 _159_ VGND 8.37f $ **FLOATING
C819 net3 VGND 3.01f $ **FLOATING
C820 a_18753_10548# VGND 0.524f $ **FLOATING
C821 ts.ts_core.dac.vdac_single.einvp_batch\[0\].pupd_47.LO VGND 0.479f $ **FLOATING
C822 net47 VGND 4.12f $ **FLOATING
C823 a_16569_10383# VGND 0.824f $ **FLOATING
C824 ts.ts_core.dac.vdac_single.en_pupd VGND 2.74f $ **FLOATING
C825 a_15315_10383# VGND 0.277f $ **FLOATING
C826 a_15125_10383# VGND 0.168f $ **FLOATING
C827 a_14857_10383# VGND 0.289f $ **FLOATING
C828 a_16591_10645# VGND 1.18f $ **FLOATING
C829 _069_ VGND 6.81f $ **FLOATING
C830 a_15959_10633# VGND 0.388f $ **FLOATING
C831 _094_ VGND 5.86f $ **FLOATING
C832 a_8856_10383# VGND 0.482f $ **FLOATING
C833 _090_ VGND 5.98f $ **FLOATING
C834 _080_ VGND 0.894f $ **FLOATING
C835 a_10516_10633# VGND 0.259f $ **FLOATING
C836 a_9687_10633# VGND 0.333f $ **FLOATING
C837 a_9290_10633# VGND 0.171f $ **FLOATING
C838 a_8938_10633# VGND 0.14f $ **FLOATING
C839 a_4883_10749# VGND 0.168f $ **FLOATING
C840 a_4680_10383# VGND 0.259f $ **FLOATING
C841 _152_ VGND 1.28f $ **FLOATING
C842 a_18109_10548# VGND 0.524f $ **FLOATING
C843 a_16403_10383# VGND 1.46f $ **FLOATING
C844 a_15535_10357# VGND 0.705f $ **FLOATING
C845 a_14015_10357# VGND 0.74f $ **FLOATING
C846 a_13905_10535# VGND 0.768f $ **FLOATING
C847 a_13546_10535# VGND 0.711f $ **FLOATING
C848 a_10686_10383# VGND 0.672f $ **FLOATING
C849 _076_ VGND 0.913f $ **FLOATING
C850 a_9770_10633# VGND 0.723f $ **FLOATING
C851 _055_ VGND 1.62f $ **FLOATING
C852 a_8468_10357# VGND 1.37f $ **FLOATING
C853 a_5340_10383# VGND 0.736f $ **FLOATING
C854 a_5515_10357# VGND 0.971f $ **FLOATING
C855 a_4775_10383# VGND 0.714f $ **FLOATING
C856 a_4993_10625# VGND 0.653f $ **FLOATING
C857 a_4425_10383# VGND 1.57f $ **FLOATING
C858 a_4259_10383# VGND 1.92f $ **FLOATING
C859 a_1585_10383# VGND 0.171f $ **FLOATING
C860 a_2659_10357# VGND 0.788f $ **FLOATING
C861 a_2401_10357# VGND 0.794f $ **FLOATING
C862 a_2305_10535# VGND 0.553f $ **FLOATING
C863 net60 VGND 0.771f $ **FLOATING
C864 a_1367_10357# VGND 0.546f $ **FLOATING
C865 a_16683_10927# VGND 1.18f $ **FLOATING
C866 a_16661_11247# VGND 0.824f $ **FLOATING
C867 a_16495_10927# VGND 1.46f $ **FLOATING
C868 _075_ VGND 6.4f $ **FLOATING
C869 a_11285_10927# VGND 0.537f $ **FLOATING
C870 a_10055_10927# VGND 0.333f $ **FLOATING
C871 a_9224_10927# VGND 0.537f $ **FLOATING
C872 a_8217_10927# VGND 0.253f $ **FLOATING
C873 a_18234_10927# VGND 1.98f $ **FLOATING
C874 a_15159_11248# VGND 0.604f $ **FLOATING
C875 a_14707_10901# VGND 0.85f $ **FLOATING
C876 a_14063_10901# VGND 0.729f $ **FLOATING
C877 a_13555_10901# VGND 0.74f $ **FLOATING
C878 a_13445_11159# VGND 0.768f $ **FLOATING
C879 a_12809_11247# VGND 0.171f $ **FLOATING
C880 _079_ VGND 1.52f $ **FLOATING
C881 a_11724_11247# VGND 0.123f $ **FLOATING
C882 a_11372_11247# VGND 0.161f $ **FLOATING
C883 _127_ VGND 1.38f $ **FLOATING
C884 a_9658_11247# VGND 0.161f $ **FLOATING
C885 a_9306_11247# VGND 0.123f $ **FLOATING
C886 _054_ VGND 1.62f $ **FLOATING
C887 a_3503_10927# VGND 0.168f $ **FLOATING
C888 a_3300_11293# VGND 0.259f $ **FLOATING
C889 a_1479_10927# VGND 0.168f $ **FLOATING
C890 a_1276_11293# VGND 0.259f $ **FLOATING
C891 a_13086_11159# VGND 0.711f $ **FLOATING
C892 _078_ VGND 0.684f $ **FLOATING
C893 ts.ts_core.o_tempdelay VGND 4.68f $ **FLOATING
C894 a_12591_11159# VGND 0.546f $ **FLOATING
C895 a_11456_11247# VGND 1.37f $ **FLOATING
C896 _052_ VGND 3.71f $ **FLOATING
C897 a_10138_10927# VGND 0.723f $ **FLOATING
C898 ts.o_res\[0\] VGND 6.98f $ **FLOATING
C899 _049_ VGND 1.13f $ **FLOATING
C900 a_8836_10901# VGND 1.37f $ **FLOATING
C901 a_8386_11247# VGND 0.55f $ **FLOATING
C902 a_6945_11225# VGND 0.607f $ **FLOATING
C903 a_6516_11159# VGND 0.59f $ **FLOATING
C904 a_5381_11225# VGND 0.607f $ **FLOATING
C905 a_4952_11159# VGND 0.59f $ **FLOATING
C906 a_3960_11305# VGND 0.736f $ **FLOATING
C907 a_4135_11231# VGND 0.971f $ **FLOATING
C908 a_3395_11305# VGND 0.714f $ **FLOATING
C909 a_3613_10901# VGND 0.653f $ **FLOATING
C910 a_3045_10933# VGND 1.57f $ **FLOATING
C911 _014_ VGND 1.36f $ **FLOATING
C912 a_2879_10933# VGND 1.92f $ **FLOATING
C913 a_1936_11305# VGND 0.736f $ **FLOATING
C914 a_2111_11231# VGND 1.13f $ **FLOATING
C915 a_1371_11305# VGND 0.714f $ **FLOATING
C916 a_1589_10901# VGND 0.653f $ **FLOATING
C917 a_1021_10933# VGND 1.57f $ **FLOATING
C918 _011_ VGND 1.15f $ **FLOATING
C919 a_855_10933# VGND 1.92f $ **FLOATING
C920 a_15649_11471# VGND 0.824f $ **FLOATING
C921 a_13832_11471# VGND 0.824f $ **FLOATING
C922 net2 VGND 4.74f $ **FLOATING
C923 a_15671_11733# VGND 1.18f $ **FLOATING
C924 a_11540_11471# VGND 0.123f $ **FLOATING
C925 a_11188_11471# VGND 0.161f $ **FLOATING
C926 a_9608_11471# VGND 0.123f $ **FLOATING
C927 a_9256_11471# VGND 0.161f $ **FLOATING
C928 a_13836_11721# VGND 1.18f $ **FLOATING
C929 a_11101_11721# VGND 0.537f $ **FLOATING
C930 a_9169_11721# VGND 0.537f $ **FLOATING
C931 _048_ VGND 1.2f $ **FLOATING
C932 ts.o_res\[16\] VGND 3.57f $ **FLOATING
C933 a_6447_11837# VGND 0.168f $ **FLOATING
C934 a_6244_11471# VGND 0.259f $ **FLOATING
C935 a_18937_11636# VGND 0.524f $ **FLOATING
C936 a_17191_11445# VGND 0.698f $ **FLOATING
C937 a_15483_11471# VGND 1.46f $ **FLOATING
C938 a_14571_11623# VGND 1.46f $ **FLOATING
C939 a_11272_11471# VGND 1.37f $ **FLOATING
C940 _053_ VGND 3.62f $ **FLOATING
C941 a_9340_11471# VGND 1.37f $ **FLOATING
C942 ts.o_res\[4\] VGND 4.54f $ **FLOATING
C943 a_8532_11721# VGND 0.502f $ **FLOATING
C944 a_6904_11471# VGND 0.736f $ **FLOATING
C945 a_7079_11445# VGND 0.971f $ **FLOATING
C946 a_6339_11471# VGND 0.714f $ **FLOATING
C947 a_6557_11713# VGND 0.653f $ **FLOATING
C948 a_5989_11471# VGND 1.57f $ **FLOATING
C949 a_5823_11471# VGND 1.92f $ **FLOATING
C950 _031_ VGND 1.54f $ **FLOATING
C951 _206_ VGND 0.956f $ **FLOATING
C952 a_5043_11636# VGND 0.524f $ **FLOATING
C953 res2_n VGND 5.43f $ **FLOATING
C954 _170_ VGND 1.3f $ **FLOATING
C955 a_2695_11721# VGND 0.238f $ **FLOATING
C956 a_1585_11721# VGND 0.238f $ **FLOATING
C957 _165_ VGND 1.13f $ **FLOATING
C958 a_4680_11445# VGND 0.648f $ **FLOATING
C959 a_4135_11445# VGND 1.2f $ **FLOATING
C960 a_16683_12015# VGND 1.18f $ **FLOATING
C961 a_14567_12015# VGND 1.18f $ **FLOATING
C962 a_16661_12335# VGND 0.824f $ **FLOATING
C963 a_16495_12015# VGND 1.46f $ **FLOATING
C964 a_14545_12335# VGND 0.824f $ **FLOATING
C965 a_14379_12015# VGND 1.46f $ **FLOATING
C966 a_11359_12015# VGND 0.388f $ **FLOATING
C967 a_9500_12015# VGND 0.537f $ **FLOATING
C968 a_7929_12015# VGND 0.206f $ **FLOATING
C969 a_7285_12015# VGND 0.206f $ **FLOATING
C970 a_9934_12335# VGND 0.161f $ **FLOATING
C971 a_9582_12335# VGND 0.123f $ **FLOATING
C972 _129_ VGND 2.09f $ **FLOATING
C973 _034_ VGND 1.16f $ **FLOATING
C974 a_3779_12015# VGND 0.168f $ **FLOATING
C975 a_3576_12381# VGND 0.259f $ **FLOATING
C976 a_1775_12015# VGND 0.238f $ **FLOATING
C977 a_16180_11989# VGND 0.648f $ **FLOATING
C978 a_13595_12336# VGND 0.641f $ **FLOATING
C979 _067_ VGND 8.88f $ **FLOATING
C980 a_13231_12247# VGND 0.673f $ **FLOATING
C981 _074_ VGND 9.2f $ **FLOATING
C982 a_12603_12247# VGND 0.658f $ **FLOATING
C983 _084_ VGND 2.58f $ **FLOATING
C984 a_12313_12234# VGND 0.524f $ **FLOATING
C985 a_11851_12247# VGND 0.619f $ **FLOATING
C986 _050_ VGND 4.85f $ **FLOATING
C987 ts.o_res\[7\] VGND 4.06f $ **FLOATING
C988 _051_ VGND 5.88f $ **FLOATING
C989 a_9112_11989# VGND 1.37f $ **FLOATING
C990 a_7847_12015# VGND 0.804f $ **FLOATING
C991 a_7203_12015# VGND 0.804f $ **FLOATING
C992 ts.ts_ctrl.temp_ctr\[7\] VGND 5.6f $ **FLOATING
C993 _209_ VGND 1.06f $ **FLOATING
C994 a_6331_12234# VGND 0.524f $ **FLOATING
C995 a_4236_12393# VGND 0.736f $ **FLOATING
C996 a_4411_12319# VGND 0.971f $ **FLOATING
C997 a_3671_12393# VGND 0.714f $ **FLOATING
C998 a_3889_11989# VGND 0.653f $ **FLOATING
C999 a_3321_12021# VGND 1.57f $ **FLOATING
C1000 a_3155_12021# VGND 1.92f $ **FLOATING
C1001 a_2375_12247# VGND 0.619f $ **FLOATING
C1002 _164_ VGND 6.05f $ **FLOATING
C1003 a_16477_12559# VGND 0.824f $ **FLOATING
C1004 a_14660_12559# VGND 0.824f $ **FLOATING
C1005 a_16499_12821# VGND 1.18f $ **FLOATING
C1006 a_9792_12559# VGND 0.123f $ **FLOATING
C1007 a_9440_12559# VGND 0.161f $ **FLOATING
C1008 a_14664_12809# VGND 1.18f $ **FLOATING
C1009 _068_ VGND 8.44f $ **FLOATING
C1010 a_12752_12809# VGND 0.259f $ **FLOATING
C1011 _103_ VGND 2.03f $ **FLOATING
C1012 _119_ VGND 2.5f $ **FLOATING
C1013 _116_ VGND 1.12f $ **FLOATING
C1014 _117_ VGND 0.752f $ **FLOATING
C1015 a_10689_12809# VGND 0.206f $ **FLOATING
C1016 a_9353_12809# VGND 0.537f $ **FLOATING
C1017 _132_ VGND 1.81f $ **FLOATING
C1018 a_8749_12809# VGND 0.214f $ **FLOATING
C1019 a_8665_12809# VGND 0.167f $ **FLOATING
C1020 a_7681_12533# VGND 0.607f $ **FLOATING
C1021 a_6669_12533# VGND 0.607f $ **FLOATING
C1022 ts.o_res\[8\] VGND 4.31f $ **FLOATING
C1023 a_3435_12559# VGND 0.211f $ **FLOATING
C1024 a_4975_12925# VGND 0.168f $ **FLOATING
C1025 a_4772_12559# VGND 0.259f $ **FLOATING
C1026 a_18836_12711# VGND 0.525f $ **FLOATING
C1027 a_16311_12559# VGND 1.46f $ **FLOATING
C1028 a_15399_12711# VGND 1.46f $ **FLOATING
C1029 a_14331_12533# VGND 0.641f $ **FLOATING
C1030 a_13967_12711# VGND 0.673f $ **FLOATING
C1031 a_13603_12533# VGND 0.698f $ **FLOATING
C1032 _077_ VGND 2.02f $ **FLOATING
C1033 _070_ VGND 6.46f $ **FLOATING
C1034 a_12321_12705# VGND 0.672f $ **FLOATING
C1035 a_11343_12809# VGND 0.702f $ **FLOATING
C1036 a_10607_12809# VGND 0.804f $ **FLOATING
C1037 ts.o_res\[2\] VGND 5.88f $ **FLOATING
C1038 _088_ VGND 5.19f $ **FLOATING
C1039 a_9524_12559# VGND 1.37f $ **FLOATING
C1040 a_8583_12559# VGND 0.972f $ **FLOATING
C1041 _131_ VGND 2.53f $ **FLOATING
C1042 a_7252_12711# VGND 0.59f $ **FLOATING
C1043 a_6240_12711# VGND 0.59f $ **FLOATING
C1044 a_5432_12559# VGND 0.736f $ **FLOATING
C1045 a_5607_12533# VGND 0.971f $ **FLOATING
C1046 a_4867_12559# VGND 0.714f $ **FLOATING
C1047 a_5085_12801# VGND 0.653f $ **FLOATING
C1048 a_4517_12559# VGND 1.57f $ **FLOATING
C1049 a_4351_12559# VGND 1.92f $ **FLOATING
C1050 _013_ VGND 1.13f $ **FLOATING
C1051 _168_ VGND 3.05f $ **FLOATING
C1052 ts.ts_ctrl.temp_ctr\[4\] VGND 8.02f $ **FLOATING
C1053 a_1479_12925# VGND 0.168f $ **FLOATING
C1054 a_1276_12559# VGND 0.259f $ **FLOATING
C1055 _169_ VGND 1.24f $ **FLOATING
C1056 a_3299_12533# VGND 0.791f $ **FLOATING
C1057 a_2695_12559# VGND 0.619f $ **FLOATING
C1058 a_1936_12559# VGND 0.736f $ **FLOATING
C1059 a_2111_12533# VGND 0.971f $ **FLOATING
C1060 a_1371_12559# VGND 0.714f $ **FLOATING
C1061 a_1589_12801# VGND 0.653f $ **FLOATING
C1062 a_1021_12559# VGND 1.57f $ **FLOATING
C1063 a_855_12559# VGND 1.92f $ **FLOATING
C1064 net38 VGND 1.48f $ **FLOATING
C1065 a_16315_13103# VGND 1.18f $ **FLOATING
C1066 ts.ts_core.dac.vdac_single.einvp_batch\[0\].vref_38.HI VGND 0.415f $ **FLOATING
C1067 a_16293_13423# VGND 0.824f $ **FLOATING
C1068 a_16127_13103# VGND 1.46f $ **FLOATING
C1069 a_15259_13423# VGND 0.46f $ **FLOATING
C1070 a_14901_13423# VGND 0.326f $ **FLOATING
C1071 _059_ VGND 12.9f $ **FLOATING
C1072 a_12946_13103# VGND 0.333f $ **FLOATING
C1073 a_11977_13103# VGND 0.206f $ **FLOATING
C1074 a_11325_13103# VGND 0.214f $ **FLOATING
C1075 a_11241_13103# VGND 0.167f $ **FLOATING
C1076 a_9629_13103# VGND 0.537f $ **FLOATING
C1077 a_9025_13103# VGND 0.214f $ **FLOATING
C1078 a_8941_13103# VGND 0.167f $ **FLOATING
C1079 a_8415_13103# VGND 0.388f $ **FLOATING
C1080 a_14471_13423# VGND 0.431f $ **FLOATING
C1081 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref VGND 2.75f $ **FLOATING
C1082 a_17935_13363# VGND 1.2f $ **FLOATING
C1083 a_14015_13077# VGND 0.74f $ **FLOATING
C1084 a_13905_13335# VGND 0.768f $ **FLOATING
C1085 _101_ VGND 0.848f $ **FLOATING
C1086 _102_ VGND 0.855f $ **FLOATING
C1087 _121_ VGND 2.71f $ **FLOATING
C1088 a_10068_13423# VGND 0.123f $ **FLOATING
C1089 a_9716_13423# VGND 0.161f $ **FLOATING
C1090 _086_ VGND 2.71f $ **FLOATING
C1091 ts.o_res\[5\] VGND 4.61f $ **FLOATING
C1092 a_7183_13103# VGND 0.168f $ **FLOATING
C1093 a_6980_13469# VGND 0.259f $ **FLOATING
C1094 _192_ VGND 3.51f $ **FLOATING
C1095 _035_ VGND 1.23f $ **FLOATING
C1096 net62 VGND 1.11f $ **FLOATING
C1097 _012_ VGND 1.6f $ **FLOATING
C1098 a_13546_13335# VGND 0.711f $ **FLOATING
C1099 a_12789_13077# VGND 0.723f $ **FLOATING
C1100 a_11895_13103# VGND 0.804f $ **FLOATING
C1101 ts.ts_ctrl.temp_ctr\[5\] VGND 7.75f $ **FLOATING
C1102 a_11159_13103# VGND 0.972f $ **FLOATING
C1103 net21 VGND 4.34f $ **FLOATING
C1104 _120_ VGND 2.72f $ **FLOATING
C1105 a_9800_13423# VGND 1.37f $ **FLOATING
C1106 _047_ VGND 5.89f $ **FLOATING
C1107 a_8859_13103# VGND 0.972f $ **FLOATING
C1108 _081_ VGND 4.44f $ **FLOATING
C1109 _085_ VGND 1.36f $ **FLOATING
C1110 a_7640_13481# VGND 0.736f $ **FLOATING
C1111 a_7815_13407# VGND 0.971f $ **FLOATING
C1112 a_7075_13481# VGND 0.714f $ **FLOATING
C1113 a_7293_13077# VGND 0.653f $ **FLOATING
C1114 a_6725_13109# VGND 1.57f $ **FLOATING
C1115 a_6559_13109# VGND 1.92f $ **FLOATING
C1116 _191_ VGND 0.806f $ **FLOATING
C1117 a_5871_13335# VGND 0.619f $ **FLOATING
C1118 a_5271_13216# VGND 0.619f $ **FLOATING
C1119 _210_ VGND 1.29f $ **FLOATING
C1120 a_5043_13322# VGND 0.524f $ **FLOATING
C1121 a_4683_13077# VGND 0.788f $ **FLOATING
C1122 a_4425_13077# VGND 0.794f $ **FLOATING
C1123 a_4329_13335# VGND 0.553f $ **FLOATING
C1124 _167_ VGND 2.55f $ **FLOATING
C1125 _166_ VGND 1.22f $ **FLOATING
C1126 a_16960_13647# VGND 0.824f $ **FLOATING
C1127 a_15465_13647# VGND 0.824f $ **FLOATING
C1128 a_16964_13897# VGND 1.18f $ **FLOATING
C1129 a_15487_13909# VGND 1.18f $ **FLOATING
C1130 _071_ VGND 5.3f $ **FLOATING
C1131 _056_ VGND 2.13f $ **FLOATING
C1132 _057_ VGND 1.27f $ **FLOATING
C1133 _118_ VGND 1.41f $ **FLOATING
C1134 a_10321_13897# VGND 0.206f $ **FLOATING
C1135 a_9889_13621# VGND 0.607f $ **FLOATING
C1136 _154_ VGND 18.4f $ **FLOATING
C1137 _032_ VGND 1.21f $ **FLOATING
C1138 a_18848_13621# VGND 0.648f $ **FLOATING
C1139 net69 VGND 17.7f $ **FLOATING
C1140 a_17699_13799# VGND 1.46f $ **FLOATING
C1141 a_15299_13647# VGND 1.46f $ **FLOATING
C1142 a_14843_13621# VGND 0.74f $ **FLOATING
C1143 a_14733_13799# VGND 0.768f $ **FLOATING
C1144 a_14374_13799# VGND 0.711f $ **FLOATING
C1145 a_12157_13799# VGND 0.502f $ **FLOATING
C1146 a_10961_13799# VGND 0.502f $ **FLOATING
C1147 a_10239_13897# VGND 0.804f $ **FLOATING
C1148 ts.ts_ctrl.temp_ctr\[6\] VGND 6.25f $ **FLOATING
C1149 _082_ VGND 4.58f $ **FLOATING
C1150 a_9460_13799# VGND 0.59f $ **FLOATING
C1151 _207_ VGND 1.04f $ **FLOATING
C1152 a_7067_13812# VGND 0.524f $ **FLOATING
C1153 a_6427_13621# VGND 0.729f $ **FLOATING
C1154 a_4513_13621# VGND 4.03f $ **FLOATING
C1155 a_3307_13799# VGND 0.56f $ **FLOATING
C1156 a_17143_14191# VGND 1.18f $ **FLOATING
C1157 a_16143_14191# VGND 0.388f $ **FLOATING
C1158 net9 VGND 18f $ **FLOATING
C1159 a_17121_14511# VGND 0.824f $ **FLOATING
C1160 a_16955_14191# VGND 1.46f $ **FLOATING
C1161 _073_ VGND 10.5f $ **FLOATING
C1162 _066_ VGND 10.9f $ **FLOATING
C1163 _072_ VGND 6.07f $ **FLOATING
C1164 _083_ VGND 5.94f $ **FLOATING
C1165 a_6067_14191# VGND 0.245f $ **FLOATING
C1166 a_2951_14191# VGND 0.168f $ **FLOATING
C1167 a_2045_14191# VGND 0.238f $ **FLOATING
C1168 a_2748_14557# VGND 0.259f $ **FLOATING
C1169 a_1677_14511# VGND 0.171f $ **FLOATING
C1170 a_18671_14451# VGND 1.2f $ **FLOATING
C1171 a_16640_14165# VGND 0.648f $ **FLOATING
C1172 a_15451_14423# VGND 0.56f $ **FLOATING
C1173 net10 VGND 7.12f $ **FLOATING
C1174 a_14857_14342# VGND 0.696f $ **FLOATING
C1175 a_14379_14191# VGND 0.788f $ **FLOATING
C1176 a_14526_14165# VGND 0.795f $ **FLOATING
C1177 a_12189_14489# VGND 0.607f $ **FLOATING
C1178 a_11760_14423# VGND 0.59f $ **FLOATING
C1179 _208_ VGND 1.02f $ **FLOATING
C1180 a_9643_14410# VGND 0.524f $ **FLOATING
C1181 a_7838_14191# VGND 4.03f $ **FLOATING
C1182 clknet_0_clk VGND 11.4f $ **FLOATING
C1183 a_4259_14557# VGND 0.729f $ **FLOATING
C1184 a_3408_14569# VGND 0.736f $ **FLOATING
C1185 a_3583_14495# VGND 1.13f $ **FLOATING
C1186 a_2843_14569# VGND 0.714f $ **FLOATING
C1187 a_3061_14165# VGND 0.653f $ **FLOATING
C1188 a_2493_14197# VGND 1.57f $ **FLOATING
C1189 _015_ VGND 1.19f $ **FLOATING
C1190 a_2327_14197# VGND 1.92f $ **FLOATING
C1191 _173_ VGND 2.22f $ **FLOATING
C1192 _175_ VGND 0.765f $ **FLOATING
C1193 a_1459_14423# VGND 0.546f $ **FLOATING
C1194 a_17029_14735# VGND 0.824f $ **FLOATING
C1195 net13 VGND 7.95f $ **FLOATING
C1196 a_17051_14997# VGND 1.18f $ **FLOATING
C1197 ts.o_res\[9\] VGND 4.49f $ **FLOATING
C1198 a_12243_15101# VGND 0.168f $ **FLOATING
C1199 a_12040_14735# VGND 0.259f $ **FLOATING
C1200 a_18847_14709# VGND 0.698f $ **FLOATING
C1201 a_16863_14735# VGND 1.46f $ **FLOATING
C1202 a_12700_14735# VGND 0.736f $ **FLOATING
C1203 a_12875_14709# VGND 0.971f $ **FLOATING
C1204 a_12135_14735# VGND 0.714f $ **FLOATING
C1205 a_12353_14977# VGND 0.653f $ **FLOATING
C1206 a_11785_14735# VGND 1.57f $ **FLOATING
C1207 a_11619_14735# VGND 1.92f $ **FLOATING
C1208 _036_ VGND 1.02f $ **FLOATING
C1209 ts.o_res\[6\] VGND 3.74f $ **FLOATING
C1210 a_9759_15101# VGND 0.168f $ **FLOATING
C1211 a_9556_14735# VGND 0.259f $ **FLOATING
C1212 a_11343_14735# VGND 0.524f $ **FLOATING
C1213 _212_ VGND 0.988f $ **FLOATING
C1214 a_10216_14735# VGND 0.736f $ **FLOATING
C1215 a_10391_14709# VGND 0.971f $ **FLOATING
C1216 a_9651_14735# VGND 0.714f $ **FLOATING
C1217 a_9869_14977# VGND 0.653f $ **FLOATING
C1218 a_9301_14735# VGND 1.57f $ **FLOATING
C1219 _033_ VGND 1.12f $ **FLOATING
C1220 a_9135_14735# VGND 1.92f $ **FLOATING
C1221 ts.ts_ctrl.state\[2\] VGND 15.7f $ **FLOATING
C1222 a_3247_14735# VGND 0.18f $ **FLOATING
C1223 a_5619_15101# VGND 0.168f $ **FLOATING
C1224 a_5416_14735# VGND 0.259f $ **FLOATING
C1225 a_8399_14735# VGND 1.2f $ **FLOATING
C1226 a_8031_14735# VGND 0.524f $ **FLOATING
C1227 a_6883_14887# VGND 0.619f $ **FLOATING
C1228 a_6076_14735# VGND 0.736f $ **FLOATING
C1229 a_6251_14709# VGND 0.971f $ **FLOATING
C1230 a_5511_14735# VGND 0.714f $ **FLOATING
C1231 a_5729_14977# VGND 0.653f $ **FLOATING
C1232 a_5161_14735# VGND 1.57f $ **FLOATING
C1233 a_4995_14735# VGND 1.92f $ **FLOATING
C1234 _176_ VGND 0.941f $ **FLOATING
C1235 a_4073_14985# VGND 0.203f $ **FLOATING
C1236 _174_ VGND 1.36f $ **FLOATING
C1237 a_1479_15101# VGND 0.168f $ **FLOATING
C1238 a_1276_14735# VGND 0.259f $ **FLOATING
C1239 a_4588_14709# VGND 0.648f $ **FLOATING
C1240 a_3944_14709# VGND 0.655f $ **FLOATING
C1241 _172_ VGND 7.11f $ **FLOATING
C1242 ts.ts_ctrl.temp_ctr\[8\] VGND 6.48f $ **FLOATING
C1243 a_1936_14735# VGND 0.736f $ **FLOATING
C1244 a_2111_14709# VGND 1.54f $ **FLOATING
C1245 a_1371_14735# VGND 0.714f $ **FLOATING
C1246 a_1589_14977# VGND 0.653f $ **FLOATING
C1247 a_1021_14735# VGND 1.57f $ **FLOATING
C1248 _016_ VGND 1.17f $ **FLOATING
C1249 a_855_14735# VGND 1.92f $ **FLOATING
C1250 a_17695_15279# VGND 1.18f $ **FLOATING
C1251 a_17673_15599# VGND 0.824f $ **FLOATING
C1252 a_17507_15279# VGND 1.46f $ **FLOATING
C1253 a_12335_15279# VGND 0.168f $ **FLOATING
C1254 a_12132_15645# VGND 0.259f $ **FLOATING
C1255 a_8563_15279# VGND 0.168f $ **FLOATING
C1256 a_8360_15645# VGND 0.259f $ **FLOATING
C1257 a_6723_15279# VGND 0.168f $ **FLOATING
C1258 a_5269_15279# VGND 0.203f $ **FLOATING
C1259 a_6520_15645# VGND 0.259f $ **FLOATING
C1260 _022_ VGND 1.21f $ **FLOATING
C1261 net64 VGND 1.22f $ **FLOATING
C1262 ts.ts_core.dac_vout_ana_ VGND 0.137p $ **FLOATING
C1263 net70 VGND 10.2f $ **FLOATING
C1264 a_12792_15657# VGND 0.736f $ **FLOATING
C1265 a_12967_15583# VGND 0.971f $ **FLOATING
C1266 a_12227_15657# VGND 0.714f $ **FLOATING
C1267 a_12445_15253# VGND 0.653f $ **FLOATING
C1268 a_11877_15285# VGND 1.57f $ **FLOATING
C1269 a_11711_15285# VGND 1.92f $ **FLOATING
C1270 a_10441_15577# VGND 0.607f $ **FLOATING
C1271 a_10012_15511# VGND 0.59f $ **FLOATING
C1272 a_9020_15657# VGND 0.736f $ **FLOATING
C1273 a_9195_15583# VGND 0.971f $ **FLOATING
C1274 a_8455_15657# VGND 0.714f $ **FLOATING
C1275 a_8673_15253# VGND 0.653f $ **FLOATING
C1276 a_8105_15285# VGND 1.57f $ **FLOATING
C1277 _042_ VGND 1.12f $ **FLOATING
C1278 a_7939_15285# VGND 1.92f $ **FLOATING
C1279 a_7180_15657# VGND 0.736f $ **FLOATING
C1280 a_7355_15583# VGND 0.971f $ **FLOATING
C1281 a_6615_15657# VGND 0.714f $ **FLOATING
C1282 a_6833_15253# VGND 0.653f $ **FLOATING
C1283 a_6265_15285# VGND 1.57f $ **FLOATING
C1284 a_6099_15285# VGND 1.92f $ **FLOATING
C1285 _187_ VGND 2.46f $ **FLOATING
C1286 _190_ VGND 1.35f $ **FLOATING
C1287 _189_ VGND 1.95f $ **FLOATING
C1288 a_5140_15253# VGND 0.655f $ **FLOATING
C1289 _178_ VGND 0.824f $ **FLOATING
C1290 _179_ VGND 0.951f $ **FLOATING
C1291 a_3663_15511# VGND 0.619f $ **FLOATING
C1292 ts.ts_ctrl.temp_ctr\[9\] VGND 11.5f $ **FLOATING
C1293 a_2751_15253# VGND 0.788f $ **FLOATING
C1294 a_2493_15253# VGND 0.794f $ **FLOATING
C1295 a_2397_15511# VGND 0.553f $ **FLOATING
C1296 net11 VGND 8.62f $ **FLOATING
C1297 _037_ VGND 1.29f $ **FLOATING
C1298 ts.o_res\[10\] VGND 4.58f $ **FLOATING
C1299 a_11753_16150# VGND 0.607f $ **FLOATING
C1300 ts.o_res\[14\] VGND 3.17f $ **FLOATING
C1301 a_10495_16189# VGND 0.168f $ **FLOATING
C1302 a_10292_15823# VGND 0.259f $ **FLOATING
C1303 a_18756_15797# VGND 0.648f $ **FLOATING
C1304 _213_ VGND 0.769f $ **FLOATING
C1305 a_12587_15988# VGND 0.524f $ **FLOATING
C1306 a_12007_16150# VGND 0.59f $ **FLOATING
C1307 a_10952_15823# VGND 0.736f $ **FLOATING
C1308 a_11127_15797# VGND 0.971f $ **FLOATING
C1309 a_10387_15823# VGND 0.714f $ **FLOATING
C1310 a_10605_16065# VGND 0.653f $ **FLOATING
C1311 a_10037_15823# VGND 1.57f $ **FLOATING
C1312 a_9871_15823# VGND 1.92f $ **FLOATING
C1313 _041_ VGND 1.02f $ **FLOATING
C1314 a_8877_15797# VGND 0.607f $ **FLOATING
C1315 ts.o_res\[15\] VGND 3.96f $ **FLOATING
C1316 ts.ts_ctrl.temp_ctr\[15\] VGND 5.26f $ **FLOATING
C1317 _218_ VGND 1.23f $ **FLOATING
C1318 net58 VGND 1.28f $ **FLOATING
C1319 ts.ts_ctrl.temp_ctr\[10\] VGND 8.24f $ **FLOATING
C1320 a_3871_16189# VGND 0.168f $ **FLOATING
C1321 a_3668_15823# VGND 0.259f $ **FLOATING
C1322 a_9595_15823# VGND 0.524f $ **FLOATING
C1323 _217_ VGND 0.988f $ **FLOATING
C1324 a_8448_15975# VGND 0.59f $ **FLOATING
C1325 a_7719_15797# VGND 0.788f $ **FLOATING
C1326 a_7461_15797# VGND 0.794f $ **FLOATING
C1327 a_7365_15975# VGND 0.553f $ **FLOATING
C1328 ts.ts_ctrl.temp_ctr\[14\] VGND 6.01f $ **FLOATING
C1329 a_6983_15797# VGND 0.788f $ **FLOATING
C1330 a_6725_15797# VGND 0.794f $ **FLOATING
C1331 a_6629_15975# VGND 0.553f $ **FLOATING
C1332 a_4328_15823# VGND 0.736f $ **FLOATING
C1333 a_4503_15797# VGND 0.971f $ **FLOATING
C1334 a_3763_15823# VGND 0.714f $ **FLOATING
C1335 net18 VGND 19.2f $ **FLOATING
C1336 a_3981_16065# VGND 0.653f $ **FLOATING
C1337 a_3413_15823# VGND 1.57f $ **FLOATING
C1338 a_3247_15823# VGND 1.92f $ **FLOATING
C1339 net12 VGND 9.1f $ **FLOATING
C1340 a_6563_16687# VGND 0.211f $ **FLOATING
C1341 _021_ VGND 1.27f $ **FLOATING
C1342 _017_ VGND 1.21f $ **FLOATING
C1343 a_18847_16341# VGND 0.698f $ **FLOATING
C1344 a_9061_16665# VGND 0.607f $ **FLOATING
C1345 a_8632_16599# VGND 0.59f $ **FLOATING
C1346 a_7159_16599# VGND 0.619f $ **FLOATING
C1347 _188_ VGND 1.43f $ **FLOATING
C1348 _186_ VGND 2.26f $ **FLOATING
C1349 net66 VGND 1.13f $ **FLOATING
C1350 a_6427_16341# VGND 0.791f $ **FLOATING
C1351 a_5179_16367# VGND 1.2f $ **FLOATING
C1352 _180_ VGND 1.21f $ **FLOATING
C1353 a_3571_16586# VGND 0.524f $ **FLOATING
C1354 a_11913_16885# VGND 0.607f $ **FLOATING
C1355 ts.o_res\[11\] VGND 7.27f $ **FLOATING
C1356 a_6880_16911# VGND 0.211f $ **FLOATING
C1357 a_4713_16911# VGND 0.171f $ **FLOATING
C1358 a_9667_17277# VGND 0.168f $ **FLOATING
C1359 a_9464_16911# VGND 0.259f $ **FLOATING
C1360 a_11484_17063# VGND 0.59f $ **FLOATING
C1361 a_10124_16911# VGND 0.736f $ **FLOATING
C1362 a_10299_16885# VGND 0.971f $ **FLOATING
C1363 a_9559_16911# VGND 0.714f $ **FLOATING
C1364 a_9777_17153# VGND 0.653f $ **FLOATING
C1365 a_9209_16911# VGND 1.57f $ **FLOATING
C1366 a_9043_16911# VGND 1.92f $ **FLOATING
C1367 _038_ VGND 1.02f $ **FLOATING
C1368 a_7387_17161# VGND 0.238f $ **FLOATING
C1369 a_5081_17161# VGND 0.238f $ **FLOATING
C1370 a_8767_16911# VGND 0.524f $ **FLOATING
C1371 _214_ VGND 0.91f $ **FLOATING
C1372 a_6690_16911# VGND 0.791f $ **FLOATING
C1373 _185_ VGND 0.745f $ **FLOATING
C1374 _114_ VGND 15.5f $ **FLOATING
C1375 _184_ VGND 2.23f $ **FLOATING
C1376 _182_ VGND 1.29f $ **FLOATING
C1377 _138_ VGND 18.7f $ **FLOATING
C1378 _137_ VGND 7.66f $ **FLOATING
C1379 _181_ VGND 0.77f $ **FLOATING
C1380 a_4495_16885# VGND 0.546f $ **FLOATING
C1381 ts.o_res\[13\] VGND 4.19f $ **FLOATING
C1382 a_11875_17455# VGND 0.168f $ **FLOATING
C1383 a_11672_17821# VGND 0.259f $ **FLOATING
C1384 ts.ts_ctrl.temp_ctr\[13\] VGND 7.84f $ **FLOATING
C1385 a_7827_17455# VGND 0.168f $ **FLOATING
C1386 a_7624_17821# VGND 0.259f $ **FLOATING
C1387 _183_ VGND 1.52f $ **FLOATING
C1388 net63 VGND 1.24f $ **FLOATING
C1389 a_4239_17455# VGND 0.168f $ **FLOATING
C1390 a_4036_17821# VGND 0.259f $ **FLOATING
C1391 a_12332_17833# VGND 0.736f $ **FLOATING
C1392 a_12507_17759# VGND 0.971f $ **FLOATING
C1393 a_11767_17833# VGND 0.714f $ **FLOATING
C1394 a_11985_17429# VGND 0.653f $ **FLOATING
C1395 a_11417_17461# VGND 1.57f $ **FLOATING
C1396 _040_ VGND 1.02f $ **FLOATING
C1397 a_11251_17461# VGND 1.92f $ **FLOATING
C1398 a_10975_17455# VGND 0.524f $ **FLOATING
C1399 _216_ VGND 1.05f $ **FLOATING
C1400 a_9871_17455# VGND 0.524f $ **FLOATING
C1401 a_8284_17833# VGND 0.736f $ **FLOATING
C1402 a_8459_17759# VGND 1.13f $ **FLOATING
C1403 a_7719_17833# VGND 0.714f $ **FLOATING
C1404 a_7937_17429# VGND 0.653f $ **FLOATING
C1405 a_7369_17461# VGND 1.57f $ **FLOATING
C1406 _020_ VGND 1.23f $ **FLOATING
C1407 a_7203_17461# VGND 1.92f $ **FLOATING
C1408 _177_ VGND 8.71f $ **FLOATING
C1409 a_6607_17687# VGND 0.619f $ **FLOATING
C1410 ts.ts_ctrl.temp_ctr\[11\] VGND 8.75f $ **FLOATING
C1411 a_6247_17429# VGND 0.788f $ **FLOATING
C1412 a_5989_17429# VGND 0.794f $ **FLOATING
C1413 a_5893_17687# VGND 0.553f $ **FLOATING
C1414 a_4696_17833# VGND 0.736f $ **FLOATING
C1415 a_4871_17759# VGND 1.54f $ **FLOATING
C1416 a_4131_17833# VGND 0.714f $ **FLOATING
C1417 net20 VGND 12.1f $ **FLOATING
C1418 a_4349_17429# VGND 0.653f $ **FLOATING
C1419 a_3781_17461# VGND 1.57f $ **FLOATING
C1420 _018_ VGND 1.31f $ **FLOATING
C1421 a_3615_17461# VGND 1.92f $ **FLOATING
C1422 clknet_2_2__leaf_clk VGND 18.1f $ **FLOATING
C1423 a_10334_18365# VGND 0.259f $ **FLOATING
C1424 a_9916_18365# VGND 0.168f $ **FLOATING
C1425 a_6999_18365# VGND 0.168f $ **FLOATING
C1426 a_6796_17999# VGND 0.259f $ **FLOATING
C1427 _039_ VGND 1.25f $ **FLOATING
C1428 a_9702_18365# VGND 0.653f $ **FLOATING
C1429 a_9771_18236# VGND 0.714f $ **FLOATING
C1430 a_9615_18141# VGND 1.92f $ **FLOATING
C1431 a_9576_18267# VGND 1.57f $ **FLOATING
C1432 a_9298_18251# VGND 0.736f $ **FLOATING
C1433 a_9095_17973# VGND 0.971f $ **FLOATING
C1434 a_7456_17999# VGND 0.736f $ **FLOATING
C1435 a_7631_17973# VGND 1.13f $ **FLOATING
C1436 a_6891_17999# VGND 0.714f $ **FLOATING
C1437 net19 VGND 18.7f $ **FLOATING
C1438 a_7109_18241# VGND 0.653f $ **FLOATING
C1439 a_6541_17999# VGND 1.57f $ **FLOATING
C1440 _019_ VGND 1.75f $ **FLOATING
C1441 a_6375_17999# VGND 1.92f $ **FLOATING
C1442 clknet_2_3__leaf_clk VGND 16.4f $ **FLOATING
C1443 tt_um_hpretl_tt06_tempsens_45.HI VGND 0.415f $ **FLOATING
C1444 tt_um_hpretl_tt06_tempsens_41.HI VGND 0.415f $ **FLOATING
C1445 tt_um_hpretl_tt06_tempsens_46.HI VGND 0.415f $ **FLOATING
C1446 _215_ VGND 1.18f $ **FLOATING
C1447 tt_um_hpretl_tt06_tempsens_51.LO VGND 0.479f $ **FLOATING
C1448 net8 VGND 10f $ **FLOATING
C1449 a_9339_18582# VGND 0.59f $ **FLOATING
C1450 ts.o_res\[12\] VGND 5.54f $ **FLOATING
C1451 ts.ts_ctrl.temp_ctr\[12\] VGND 7.75f $ **FLOATING
C1452 a_9085_18582# VGND 0.607f $ **FLOATING
C1453 _211_ VGND 20.4f $ **FLOATING
C1454 a_8399_18543# VGND 1.2f $ **FLOATING
C1455 tt_um_hpretl_tt06_tempsens_48.LO VGND 0.479f $ **FLOATING
.ends
