magic
tech sky130A
magscale 1 2
timestamp 1712951395
<< nwell >>
rect 5996 -516 6090 -472
rect 5996 -518 6078 -516
rect 6062 -580 6080 -560
rect 6922 -620 6934 -616
rect 6950 -926 6984 -820
rect 7866 -900 7900 -836
<< pwell >>
rect 4878 -2100 6912 -2054
rect 4468 -2334 4514 -2286
rect 4878 -2406 6912 -2368
rect 4878 -2414 4884 -2406
rect 15972 -2516 16000 -2458
<< viali >>
rect 1928 -444 2078 -386
rect 6016 -512 8834 -478
rect 9420 -502 12238 -468
rect 16058 -984 16092 -610
rect 1908 -2088 2088 -1990
rect 5082 -2508 6984 -2474
rect 12708 -2504 15984 -2470
rect 2656 -2692 4558 -2658
rect 7574 -2694 7802 -2660
rect 10860 -2696 11084 -2626
<< metal1 >>
rect 12834 612 16136 620
rect 1516 140 16136 612
rect 1516 50 9836 140
rect 1516 40 8284 50
rect 1516 34 7364 40
rect 1516 -82 6450 34
rect 6562 -82 7364 34
rect 1516 -84 7364 -82
rect 7478 -82 8284 40
rect 8398 -62 9836 50
rect 9986 138 16136 140
rect 9986 134 11658 138
rect 9986 -62 10752 134
rect 8398 -68 10752 -62
rect 10902 -64 11658 134
rect 11808 112 16136 138
rect 11808 -64 12948 112
rect 10902 -68 12948 -64
rect 8398 -78 12948 -68
rect 15694 -78 16136 112
rect 8398 -82 16136 -78
rect 7478 -84 16136 -82
rect 1516 -86 16136 -84
rect 1516 -88 2772 -86
rect 1522 -246 1718 -240
rect 1522 -386 2246 -246
rect 1522 -444 1928 -386
rect 2078 -444 2246 -386
rect 1522 -452 2246 -444
rect 1522 -2804 1718 -452
rect 2340 -482 2772 -88
rect 6016 -466 8834 -86
rect 9422 -394 16136 -86
rect 9422 -446 12240 -394
rect 9408 -450 12240 -446
rect 1798 -914 2772 -482
rect 5996 -478 8850 -466
rect 5996 -512 6016 -478
rect 8834 -512 8850 -478
rect 9408 -468 12262 -450
rect 9408 -502 9420 -468
rect 12238 -502 12262 -468
rect 12758 -488 16136 -394
rect 9408 -508 12262 -502
rect 5996 -518 8850 -512
rect 12174 -514 12262 -508
rect 12738 -526 16136 -488
rect 16018 -560 16136 -526
rect 5320 -580 5868 -562
rect 6084 -580 6476 -574
rect 9484 -580 9884 -564
rect 9946 -580 10796 -564
rect 10860 -580 11254 -564
rect 11316 -580 11710 -564
rect 11774 -580 12168 -564
rect 5320 -616 8722 -580
rect 8738 -614 12173 -580
rect 16032 -610 16136 -560
rect 5320 -896 5838 -616
rect 6008 -672 6046 -616
rect 6084 -620 6476 -616
rect 6542 -620 6934 -616
rect 6008 -840 6068 -672
rect 6008 -856 6072 -840
rect 6438 -856 6448 -658
rect 6562 -856 6572 -658
rect 6950 -670 6984 -648
rect 6950 -848 6986 -670
rect 6008 -896 6046 -856
rect 6950 -896 6984 -848
rect 7356 -862 7366 -664
rect 7480 -862 7490 -664
rect 7866 -846 7902 -676
rect 7866 -896 7900 -846
rect 8272 -862 8282 -664
rect 8396 -862 8406 -664
rect 8780 -896 8814 -672
rect 9018 -896 9254 -614
rect 12468 -616 12670 -610
rect 12834 -616 12926 -610
rect 13000 -616 15929 -610
rect 12468 -644 15929 -616
rect 12132 -646 15929 -644
rect 9372 -852 9382 -650
rect 9532 -852 9542 -650
rect 9830 -854 9840 -652
rect 9990 -854 10000 -652
rect 10280 -852 10290 -650
rect 10440 -852 10450 -650
rect 10742 -850 10752 -648
rect 10902 -850 10912 -648
rect 11198 -854 11208 -652
rect 11358 -854 11368 -652
rect 11656 -854 11666 -652
rect 11816 -854 11826 -652
rect 12120 -848 12130 -646
rect 12280 -656 15929 -646
rect 12280 -848 12714 -656
rect 12132 -852 12714 -848
rect 1798 -1112 2230 -914
rect 5320 -942 12172 -896
rect 5322 -948 12172 -942
rect 12468 -938 12714 -852
rect 12764 -896 12774 -690
rect 12830 -896 12840 -690
rect 12920 -904 12930 -698
rect 12986 -904 12996 -698
rect 13080 -902 13090 -696
rect 13146 -902 13156 -696
rect 13234 -900 13244 -694
rect 13300 -900 13310 -694
rect 13392 -902 13402 -696
rect 13458 -902 13468 -696
rect 13550 -902 13560 -696
rect 13616 -902 13626 -696
rect 13712 -900 13722 -694
rect 13778 -900 13788 -694
rect 13868 -902 13878 -696
rect 13934 -902 13944 -696
rect 14028 -900 14038 -694
rect 14094 -900 14104 -694
rect 14186 -900 14196 -694
rect 14252 -900 14262 -694
rect 14342 -902 14352 -696
rect 14408 -902 14418 -696
rect 14500 -902 14510 -696
rect 14566 -902 14576 -696
rect 14658 -900 14668 -694
rect 14724 -900 14734 -694
rect 14816 -902 14826 -696
rect 14882 -902 14892 -696
rect 14972 -902 14982 -696
rect 15038 -902 15048 -696
rect 15130 -902 15140 -696
rect 15196 -902 15206 -696
rect 15288 -902 15298 -696
rect 15354 -902 15364 -696
rect 15450 -898 15460 -692
rect 15516 -898 15526 -692
rect 15606 -898 15616 -692
rect 15672 -898 15682 -692
rect 15762 -902 15772 -696
rect 15828 -902 15838 -696
rect 15922 -904 15932 -698
rect 15988 -904 15998 -698
rect 5322 -950 5838 -948
rect 7710 -1062 8696 -948
rect 12468 -984 15929 -938
rect 16032 -984 16058 -610
rect 16092 -984 16136 -610
rect 7972 -1140 8116 -1062
rect 16032 -1110 16136 -984
rect 4506 -1362 7873 -1243
rect 7962 -1280 7972 -1140
rect 8112 -1280 8122 -1140
rect 13146 -1258 15844 -1230
rect 4506 -1492 12463 -1362
rect 4480 -1494 12463 -1492
rect 1782 -1665 12463 -1494
rect 13146 -1466 13176 -1258
rect 15788 -1378 15844 -1258
rect 15788 -1398 15936 -1378
rect 15788 -1466 16084 -1398
rect 13146 -1568 16084 -1466
rect 15704 -1598 16084 -1568
rect 15704 -1628 16022 -1598
rect 1782 -1914 4930 -1665
rect 7452 -1680 12463 -1665
rect 15862 -1670 16022 -1628
rect 7452 -1712 12464 -1680
rect 1788 -1990 2212 -1974
rect 1788 -2088 1908 -1990
rect 2088 -2088 2212 -1990
rect 1788 -2804 2212 -2088
rect 2316 -2314 2524 -1914
rect 2736 -2280 3104 -1914
rect 3194 -2080 3570 -1914
rect 3194 -2280 3564 -2080
rect 3652 -2280 4020 -1914
rect 4110 -2206 4478 -1914
rect 4836 -2054 4930 -1914
rect 7174 -1894 9639 -1752
rect 4836 -2100 6912 -2054
rect 4110 -2280 4480 -2206
rect 2316 -2522 2726 -2314
rect 3048 -2514 3058 -2318
rect 3228 -2514 3238 -2318
rect 3278 -2320 3460 -2280
rect 3746 -2320 3928 -2280
rect 4278 -2286 4480 -2280
rect 3278 -2514 3938 -2320
rect 3974 -2514 3984 -2318
rect 4154 -2514 4164 -2318
rect 4278 -2328 4514 -2286
rect 4278 -2514 4548 -2328
rect 4836 -2368 4930 -2100
rect 5024 -2326 5034 -2142
rect 5220 -2326 5230 -2142
rect 5434 -2330 5444 -2132
rect 5702 -2330 5712 -2132
rect 5936 -2322 5946 -2138
rect 6132 -2322 6142 -2138
rect 6350 -2334 6360 -2136
rect 6618 -2334 6628 -2136
rect 6850 -2328 6860 -2144
rect 7046 -2146 7056 -2144
rect 7174 -2146 7316 -1894
rect 7638 -1982 8400 -1948
rect 7046 -2324 7626 -2146
rect 7750 -2168 8166 -2030
rect 7750 -2324 7972 -2168
rect 8112 -2324 8166 -2168
rect 7046 -2328 7056 -2324
rect 4836 -2406 6912 -2368
rect 4836 -2414 4884 -2406
rect 4944 -2470 7106 -2468
rect 4944 -2474 7112 -2470
rect 4944 -2508 5082 -2474
rect 6984 -2508 7112 -2474
rect 7750 -2508 8166 -2324
rect 8366 -2414 8400 -1982
rect 9497 -2147 9639 -1894
rect 10065 -1947 11027 -1909
rect 9491 -2289 9497 -2147
rect 9639 -2289 9645 -2147
rect 10065 -2410 10103 -1947
rect 10215 -2150 10922 -2120
rect 10205 -2289 10215 -2150
rect 10586 -2289 10922 -2150
rect 11032 -2156 11600 -1986
rect 3278 -2516 3460 -2514
rect 3746 -2518 3928 -2514
rect 2316 -2524 2524 -2522
rect 2316 -2552 2442 -2524
rect 2316 -2590 4512 -2552
rect 4944 -2578 7112 -2508
rect 8328 -2558 8528 -2414
rect 2316 -2648 2442 -2590
rect 2560 -2654 4708 -2652
rect 2560 -2658 4712 -2654
rect 2560 -2692 2656 -2658
rect 4558 -2692 4712 -2658
rect 2560 -2758 4712 -2692
rect 2560 -2804 3060 -2758
rect 1522 -2918 3060 -2804
rect 3230 -2918 3986 -2758
rect 4156 -2804 4712 -2758
rect 4944 -2804 5438 -2578
rect 4156 -2816 5438 -2804
rect 6634 -2804 7112 -2578
rect 7636 -2592 8528 -2558
rect 8328 -2614 8528 -2592
rect 9870 -2518 10103 -2410
rect 11032 -2388 11424 -2156
rect 11566 -2388 11600 -2156
rect 11032 -2478 11600 -2388
rect 12106 -2056 12464 -1712
rect 13152 -1710 16022 -1670
rect 13152 -1882 13184 -1710
rect 15938 -1882 16022 -1710
rect 13152 -1904 16022 -1882
rect 12106 -2098 15928 -2056
rect 12106 -2362 12464 -2098
rect 12690 -2326 12700 -2126
rect 12782 -2326 12792 -2126
rect 13146 -2328 13156 -2128
rect 13238 -2328 13248 -2128
rect 13606 -2326 13616 -2126
rect 13698 -2326 13708 -2126
rect 14072 -2332 14082 -2132
rect 14164 -2332 14174 -2132
rect 14522 -2326 14532 -2126
rect 14614 -2326 14624 -2126
rect 14980 -2328 14990 -2128
rect 15072 -2328 15082 -2128
rect 15440 -2328 15450 -2128
rect 15532 -2328 15542 -2128
rect 15898 -2332 15908 -2132
rect 15990 -2332 16000 -2132
rect 12106 -2404 15922 -2362
rect 12106 -2418 12464 -2404
rect 12696 -2464 12724 -2458
rect 15972 -2464 16000 -2458
rect 12696 -2470 16000 -2464
rect 12696 -2504 12708 -2470
rect 15984 -2504 16000 -2470
rect 12696 -2516 16000 -2504
rect 9870 -2556 11022 -2518
rect 9870 -2610 10070 -2556
rect 10854 -2624 11090 -2618
rect 10736 -2626 11186 -2624
rect 7464 -2660 7912 -2646
rect 7464 -2694 7574 -2660
rect 7802 -2694 7912 -2660
rect 7464 -2804 7912 -2694
rect 10736 -2696 10860 -2626
rect 11084 -2696 11186 -2626
rect 10736 -2804 11186 -2696
rect 12706 -2804 15990 -2516
rect 6634 -2816 16105 -2804
rect 4156 -2844 16105 -2816
rect 4156 -2918 12694 -2844
rect 1522 -3032 12694 -2918
rect 16002 -3032 16105 -2844
rect 1522 -3502 16105 -3032
rect 1522 -3504 1718 -3502
<< via1 >>
rect 6450 -82 6562 34
rect 7364 -84 7478 40
rect 8284 -82 8398 50
rect 9836 -62 9986 140
rect 10752 -68 10902 134
rect 11658 -64 11808 138
rect 12948 -78 15694 112
rect 6448 -856 6562 -658
rect 7366 -862 7480 -664
rect 8282 -862 8396 -664
rect 9382 -852 9532 -650
rect 9840 -854 9990 -652
rect 10290 -852 10440 -650
rect 10752 -850 10902 -648
rect 11208 -854 11358 -652
rect 11666 -854 11816 -652
rect 12130 -848 12280 -646
rect 12774 -896 12830 -690
rect 12930 -904 12986 -698
rect 13090 -902 13146 -696
rect 13244 -900 13300 -694
rect 13402 -902 13458 -696
rect 13560 -902 13616 -696
rect 13722 -900 13778 -694
rect 13878 -902 13934 -696
rect 14038 -900 14094 -694
rect 14196 -900 14252 -694
rect 14352 -902 14408 -696
rect 14510 -902 14566 -696
rect 14668 -900 14724 -694
rect 14826 -902 14882 -696
rect 14982 -902 15038 -696
rect 15140 -902 15196 -696
rect 15298 -902 15354 -696
rect 15460 -898 15516 -692
rect 15616 -898 15672 -692
rect 15772 -902 15828 -696
rect 15932 -904 15988 -698
rect 7972 -1280 8112 -1140
rect 13176 -1466 15788 -1258
rect 3058 -2514 3228 -2318
rect 3984 -2514 4154 -2318
rect 5034 -2326 5220 -2142
rect 5444 -2330 5702 -2132
rect 5946 -2322 6132 -2138
rect 6360 -2334 6618 -2136
rect 6860 -2328 7046 -2144
rect 7972 -2324 8112 -2168
rect 9497 -2289 9639 -2147
rect 10215 -2289 10586 -2150
rect 3060 -2918 3230 -2758
rect 3986 -2918 4156 -2758
rect 5438 -2816 6634 -2578
rect 11424 -2388 11566 -2156
rect 13184 -1882 15938 -1710
rect 12700 -2326 12782 -2126
rect 13156 -2328 13238 -2128
rect 13616 -2326 13698 -2126
rect 14082 -2332 14164 -2132
rect 14532 -2326 14614 -2126
rect 14990 -2328 15072 -2128
rect 15450 -2328 15532 -2128
rect 15908 -2332 15990 -2132
rect 12694 -3032 16002 -2844
<< metal2 >>
rect 9836 140 9986 150
rect 8284 50 8398 60
rect 6450 36 6562 44
rect 6448 34 6562 36
rect 6448 -82 6450 34
rect 6448 -658 6562 -82
rect 7364 40 7478 50
rect 7478 -84 7482 -8
rect 7364 -94 7482 -84
rect 6438 -856 6448 -658
rect 6562 -856 6572 -658
rect 7366 -664 7482 -94
rect 9836 -72 9986 -62
rect 10752 134 10902 144
rect 8284 -92 8398 -82
rect 8284 -654 8394 -92
rect 9382 -644 9532 -640
rect 9848 -642 9982 -72
rect 10752 -78 10902 -68
rect 11658 138 11808 148
rect 11658 -74 11808 -64
rect 12926 112 15842 128
rect 10756 -638 10890 -78
rect 9382 -650 9536 -644
rect 8284 -664 8396 -654
rect 6448 -866 6562 -856
rect 7356 -862 7366 -664
rect 7480 -862 7490 -664
rect 8272 -862 8282 -664
rect 8396 -862 8406 -664
rect 9532 -852 9536 -650
rect 9382 -862 9536 -852
rect 7366 -872 7480 -862
rect 8282 -872 8396 -862
rect 9384 -998 9536 -862
rect 9840 -652 9990 -642
rect 9840 -864 9990 -854
rect 10290 -650 10440 -640
rect 10290 -862 10440 -852
rect 10752 -648 10902 -638
rect 11670 -642 11804 -74
rect 12926 -78 12948 112
rect 15694 -78 15842 112
rect 12926 -426 15842 -78
rect 10752 -860 10902 -850
rect 11208 -652 11358 -642
rect 10292 -998 10432 -862
rect 11208 -864 11358 -854
rect 11666 -652 11816 -642
rect 11666 -862 11816 -854
rect 12130 -646 12280 -636
rect 12130 -858 12280 -848
rect 12766 -690 12832 -680
rect 11212 -998 11352 -864
rect 12130 -998 12270 -858
rect 7972 -1140 8112 -1130
rect 9384 -1188 12270 -998
rect 12766 -896 12774 -690
rect 12830 -896 12832 -690
rect 12766 -1170 12832 -896
rect 12926 -698 12992 -426
rect 12926 -904 12930 -698
rect 12986 -904 12992 -698
rect 12926 -914 12992 -904
rect 13084 -696 13150 -686
rect 13084 -902 13090 -696
rect 13146 -902 13150 -696
rect 13084 -1170 13150 -902
rect 13240 -694 13306 -426
rect 13402 -690 13458 -686
rect 13240 -900 13244 -694
rect 13300 -900 13306 -694
rect 13240 -906 13306 -900
rect 13398 -696 13464 -690
rect 13398 -902 13402 -696
rect 13458 -902 13464 -696
rect 13244 -910 13300 -906
rect 13398 -1170 13464 -902
rect 13554 -696 13620 -426
rect 13554 -902 13560 -696
rect 13616 -902 13620 -696
rect 13554 -906 13620 -902
rect 13718 -694 13784 -684
rect 13718 -900 13722 -694
rect 13778 -900 13784 -694
rect 13560 -912 13616 -906
rect 13718 -1170 13784 -900
rect 13872 -696 13938 -426
rect 13872 -902 13878 -696
rect 13934 -902 13938 -696
rect 13872 -916 13938 -902
rect 14032 -694 14098 -684
rect 14032 -900 14038 -694
rect 14094 -900 14098 -694
rect 14032 -1170 14098 -900
rect 14192 -694 14258 -426
rect 14352 -688 14408 -686
rect 14192 -900 14196 -694
rect 14252 -900 14258 -694
rect 14192 -904 14258 -900
rect 14346 -696 14412 -688
rect 14346 -902 14352 -696
rect 14408 -902 14412 -696
rect 14196 -910 14252 -904
rect 14346 -1170 14412 -902
rect 14504 -696 14570 -426
rect 14504 -902 14510 -696
rect 14566 -902 14570 -696
rect 14504 -906 14570 -902
rect 14660 -694 14726 -684
rect 14660 -900 14668 -694
rect 14724 -900 14726 -694
rect 14510 -912 14566 -906
rect 14660 -1170 14726 -900
rect 14822 -696 14888 -426
rect 14982 -692 15038 -686
rect 14822 -902 14826 -696
rect 14882 -902 14888 -696
rect 14822 -908 14888 -902
rect 14976 -696 15042 -692
rect 14976 -902 14982 -696
rect 15038 -902 15042 -696
rect 14826 -912 14882 -908
rect 14976 -1170 15042 -902
rect 15136 -696 15202 -426
rect 15298 -688 15354 -686
rect 15136 -902 15140 -696
rect 15196 -902 15202 -696
rect 15136 -906 15202 -902
rect 15296 -696 15362 -688
rect 15296 -902 15298 -696
rect 15354 -902 15362 -696
rect 15140 -912 15196 -906
rect 15296 -1170 15362 -902
rect 15454 -692 15520 -426
rect 15616 -692 15672 -682
rect 15454 -898 15460 -692
rect 15516 -898 15520 -692
rect 15454 -906 15520 -898
rect 15610 -898 15616 -692
rect 15672 -898 15676 -692
rect 15460 -908 15516 -906
rect 15610 -1170 15676 -898
rect 15766 -696 15832 -426
rect 15766 -902 15772 -696
rect 15828 -902 15832 -696
rect 15766 -904 15832 -902
rect 15928 -698 15994 -686
rect 15928 -904 15932 -698
rect 15988 -904 15994 -698
rect 15772 -912 15828 -904
rect 15928 -1170 15994 -904
rect 5034 -1966 7045 -1776
rect 5034 -2142 5224 -1966
rect 3058 -2312 3228 -2308
rect 3058 -2318 3230 -2312
rect 3228 -2514 3230 -2318
rect 3058 -2758 3230 -2514
rect 3984 -2318 4156 -2308
rect 4154 -2514 4156 -2318
rect 5220 -2326 5224 -2142
rect 5444 -2130 5702 -2122
rect 5947 -2128 6137 -1966
rect 5444 -2132 5708 -2130
rect 5034 -2336 5220 -2326
rect 5702 -2330 5708 -2132
rect 3984 -2524 4156 -2514
rect 3988 -2748 4156 -2524
rect 5444 -2568 5708 -2330
rect 5946 -2138 6137 -2128
rect 6132 -2322 6137 -2138
rect 5946 -2325 6137 -2322
rect 6360 -2128 6618 -2126
rect 6360 -2136 6628 -2128
rect 5946 -2332 6132 -2325
rect 6618 -2334 6628 -2136
rect 6855 -2134 7045 -1966
rect 6855 -2144 7046 -2134
rect 6855 -2328 6860 -2144
rect 6855 -2333 7046 -2328
rect 6360 -2344 6628 -2334
rect 6860 -2338 7046 -2333
rect 7972 -2168 8112 -1280
rect 11424 -1190 12270 -1188
rect 9497 -2147 9639 -2141
rect 10215 -2147 10586 -2140
rect 9639 -2150 10586 -2147
rect 9639 -2289 10215 -2150
rect 9497 -2295 9639 -2289
rect 10215 -2299 10586 -2289
rect 11424 -2156 11576 -1190
rect 12744 -1214 16094 -1170
rect 12740 -1258 16094 -1214
rect 12740 -1466 13176 -1258
rect 15788 -1342 16094 -1258
rect 15788 -1466 15824 -1342
rect 12740 -1480 15824 -1466
rect 13184 -1708 15938 -1700
rect 13164 -1710 16000 -1708
rect 13164 -1814 13184 -1710
rect 13160 -1882 13184 -1814
rect 15938 -1882 16000 -1710
rect 13160 -1896 16000 -1882
rect 7972 -2334 8112 -2324
rect 6364 -2568 6628 -2344
rect 11566 -2386 11576 -2156
rect 12700 -2126 12782 -2116
rect 13160 -2118 13236 -1896
rect 12700 -2336 12782 -2326
rect 13156 -2128 13238 -2118
rect 11424 -2398 11566 -2388
rect 3058 -2918 3060 -2758
rect 3058 -2920 3230 -2918
rect 3060 -2928 3230 -2920
rect 3986 -2758 4156 -2748
rect 5438 -2578 6634 -2568
rect 5438 -2826 6634 -2816
rect 12700 -2834 12776 -2336
rect 13156 -2338 13238 -2328
rect 13616 -2126 13698 -2116
rect 13616 -2336 13698 -2326
rect 14080 -2122 14156 -1896
rect 14080 -2132 14164 -2122
rect 14080 -2332 14082 -2132
rect 14080 -2336 14164 -2332
rect 14532 -2126 14614 -2116
rect 14532 -2336 14614 -2326
rect 13620 -2834 13696 -2336
rect 14082 -2342 14164 -2336
rect 14538 -2834 14614 -2336
rect 14990 -2118 15066 -1896
rect 14990 -2128 15072 -2118
rect 14990 -2338 15072 -2328
rect 15450 -2128 15532 -2118
rect 15912 -2122 15988 -1896
rect 15450 -2338 15532 -2328
rect 15908 -2132 15990 -2122
rect 15454 -2834 15530 -2338
rect 15908 -2342 15990 -2332
rect 3986 -2928 4156 -2918
rect 12694 -2844 16002 -2834
rect 12694 -3042 16002 -3032
use sky130_fd_pr__nfet_01v8_lvt_8TELWR  XM1
timestamp 1712811291
transform 1 0 10972 0 1 -2234
box -246 -460 246 460
use sky130_fd_pr__nfet_01v8_lvt_8TELWR  XM2
timestamp 1712811291
transform 1 0 7688 0 1 -2270
box -246 -460 246 460
use sky130_fd_pr__nfet_01v8_VWWVRL  XM3
timestamp 1712811291
transform 1 0 6033 0 1 -2234
box -1083 -310 1083 310
use sky130_fd_pr__pfet_01v8_lvt_GW6ZVV  XM4
timestamp 1712811291
transform 1 0 7425 0 1 -761
box -1541 -319 1541 319
use sky130_fd_pr__pfet_01v8_lvt_GW6ZVV  XM5
timestamp 1712811291
transform 1 0 10829 0 1 -751
box -1541 -319 1541 319
use sky130_fd_pr__nfet_01v8_VWWVRL  XM6
timestamp 1712811291
transform 1 0 3607 0 1 -2418
box -1083 -310 1083 310
use sky130_fd_pr__nfet_01v8_WWWVRA  XM7
timestamp 1712811291
transform 1 0 14346 0 1 -2230
box -1770 -310 1770 310
use sky130_fd_pr__pfet_01v8_lvt_ER3WAW  XM8
timestamp 1712811291
transform 1 0 14381 0 1 -797
box -1747 -319 1747 319
use sky130_fd_pr__res_xhigh_po_0p35_5BGKUX  XR1
timestamp 1712811291
transform 1 0 2005 0 1 -1232
box -201 -862 201 862
<< labels >>
flabel metal1 1806 314 2006 514 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1800 -3080 2000 -2880 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 8328 -2614 8528 -2414 0 FreeSans 256 0 0 0 MINUS
port 1 nsew
flabel metal1 9870 -2610 10070 -2410 0 FreeSans 256 0 0 0 PLUS
port 2 nsew
flabel metal1 15884 -1598 16084 -1398 0 FreeSans 256 0 0 0 VOUT
port 3 nsew
flabel metal1 1782 -1914 4930 -1494 0 FreeSans 480 0 0 0 VBIAS
flabel metal1 9497 -2147 9639 -1752 0 FreeSans 480 0 0 0 VX
flabel space 7744 -2508 8166 -2324 0 FreeSans 480 0 0 0 V2
flabel space 11028 -2478 11424 -1986 0 FreeSans 480 0 0 0 V1
<< end >>
