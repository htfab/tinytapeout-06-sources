magic
tech sky130A
timestamp 1713448216
<< pwell >>
rect -148 -8368 148 8368
<< nmos >>
rect -50 7263 50 8263
rect -50 6154 50 7154
rect -50 5045 50 6045
rect -50 3936 50 4936
rect -50 2827 50 3827
rect -50 1718 50 2718
rect -50 609 50 1609
rect -50 -500 50 500
rect -50 -1609 50 -609
rect -50 -2718 50 -1718
rect -50 -3827 50 -2827
rect -50 -4936 50 -3936
rect -50 -6045 50 -5045
rect -50 -7154 50 -6154
rect -50 -8263 50 -7263
<< ndiff >>
rect -79 8257 -50 8263
rect -79 7269 -73 8257
rect -56 7269 -50 8257
rect -79 7263 -50 7269
rect 50 8257 79 8263
rect 50 7269 56 8257
rect 73 7269 79 8257
rect 50 7263 79 7269
rect -79 7148 -50 7154
rect -79 6160 -73 7148
rect -56 6160 -50 7148
rect -79 6154 -50 6160
rect 50 7148 79 7154
rect 50 6160 56 7148
rect 73 6160 79 7148
rect 50 6154 79 6160
rect -79 6039 -50 6045
rect -79 5051 -73 6039
rect -56 5051 -50 6039
rect -79 5045 -50 5051
rect 50 6039 79 6045
rect 50 5051 56 6039
rect 73 5051 79 6039
rect 50 5045 79 5051
rect -79 4930 -50 4936
rect -79 3942 -73 4930
rect -56 3942 -50 4930
rect -79 3936 -50 3942
rect 50 4930 79 4936
rect 50 3942 56 4930
rect 73 3942 79 4930
rect 50 3936 79 3942
rect -79 3821 -50 3827
rect -79 2833 -73 3821
rect -56 2833 -50 3821
rect -79 2827 -50 2833
rect 50 3821 79 3827
rect 50 2833 56 3821
rect 73 2833 79 3821
rect 50 2827 79 2833
rect -79 2712 -50 2718
rect -79 1724 -73 2712
rect -56 1724 -50 2712
rect -79 1718 -50 1724
rect 50 2712 79 2718
rect 50 1724 56 2712
rect 73 1724 79 2712
rect 50 1718 79 1724
rect -79 1603 -50 1609
rect -79 615 -73 1603
rect -56 615 -50 1603
rect -79 609 -50 615
rect 50 1603 79 1609
rect 50 615 56 1603
rect 73 615 79 1603
rect 50 609 79 615
rect -79 494 -50 500
rect -79 -494 -73 494
rect -56 -494 -50 494
rect -79 -500 -50 -494
rect 50 494 79 500
rect 50 -494 56 494
rect 73 -494 79 494
rect 50 -500 79 -494
rect -79 -615 -50 -609
rect -79 -1603 -73 -615
rect -56 -1603 -50 -615
rect -79 -1609 -50 -1603
rect 50 -615 79 -609
rect 50 -1603 56 -615
rect 73 -1603 79 -615
rect 50 -1609 79 -1603
rect -79 -1724 -50 -1718
rect -79 -2712 -73 -1724
rect -56 -2712 -50 -1724
rect -79 -2718 -50 -2712
rect 50 -1724 79 -1718
rect 50 -2712 56 -1724
rect 73 -2712 79 -1724
rect 50 -2718 79 -2712
rect -79 -2833 -50 -2827
rect -79 -3821 -73 -2833
rect -56 -3821 -50 -2833
rect -79 -3827 -50 -3821
rect 50 -2833 79 -2827
rect 50 -3821 56 -2833
rect 73 -3821 79 -2833
rect 50 -3827 79 -3821
rect -79 -3942 -50 -3936
rect -79 -4930 -73 -3942
rect -56 -4930 -50 -3942
rect -79 -4936 -50 -4930
rect 50 -3942 79 -3936
rect 50 -4930 56 -3942
rect 73 -4930 79 -3942
rect 50 -4936 79 -4930
rect -79 -5051 -50 -5045
rect -79 -6039 -73 -5051
rect -56 -6039 -50 -5051
rect -79 -6045 -50 -6039
rect 50 -5051 79 -5045
rect 50 -6039 56 -5051
rect 73 -6039 79 -5051
rect 50 -6045 79 -6039
rect -79 -6160 -50 -6154
rect -79 -7148 -73 -6160
rect -56 -7148 -50 -6160
rect -79 -7154 -50 -7148
rect 50 -6160 79 -6154
rect 50 -7148 56 -6160
rect 73 -7148 79 -6160
rect 50 -7154 79 -7148
rect -79 -7269 -50 -7263
rect -79 -8257 -73 -7269
rect -56 -8257 -50 -7269
rect -79 -8263 -50 -8257
rect 50 -7269 79 -7263
rect 50 -8257 56 -7269
rect 73 -8257 79 -7269
rect 50 -8263 79 -8257
<< ndiffc >>
rect -73 7269 -56 8257
rect 56 7269 73 8257
rect -73 6160 -56 7148
rect 56 6160 73 7148
rect -73 5051 -56 6039
rect 56 5051 73 6039
rect -73 3942 -56 4930
rect 56 3942 73 4930
rect -73 2833 -56 3821
rect 56 2833 73 3821
rect -73 1724 -56 2712
rect 56 1724 73 2712
rect -73 615 -56 1603
rect 56 615 73 1603
rect -73 -494 -56 494
rect 56 -494 73 494
rect -73 -1603 -56 -615
rect 56 -1603 73 -615
rect -73 -2712 -56 -1724
rect 56 -2712 73 -1724
rect -73 -3821 -56 -2833
rect 56 -3821 73 -2833
rect -73 -4930 -56 -3942
rect 56 -4930 73 -3942
rect -73 -6039 -56 -5051
rect 56 -6039 73 -5051
rect -73 -7148 -56 -6160
rect 56 -7148 73 -6160
rect -73 -8257 -56 -7269
rect 56 -8257 73 -7269
<< psubdiff >>
rect -130 8333 -82 8350
rect 82 8333 130 8350
rect -130 8302 -113 8333
rect 113 8302 130 8333
rect -130 -8333 -113 -8302
rect 113 -8333 130 -8302
rect -130 -8350 -82 -8333
rect 82 -8350 130 -8333
<< psubdiffcont >>
rect -82 8333 82 8350
rect -130 -8302 -113 8302
rect 113 -8302 130 8302
rect -82 -8350 82 -8333
<< poly >>
rect -50 8299 50 8307
rect -50 8282 -42 8299
rect 42 8282 50 8299
rect -50 8263 50 8282
rect -50 7244 50 7263
rect -50 7227 -42 7244
rect 42 7227 50 7244
rect -50 7219 50 7227
rect -50 7190 50 7198
rect -50 7173 -42 7190
rect 42 7173 50 7190
rect -50 7154 50 7173
rect -50 6135 50 6154
rect -50 6118 -42 6135
rect 42 6118 50 6135
rect -50 6110 50 6118
rect -50 6081 50 6089
rect -50 6064 -42 6081
rect 42 6064 50 6081
rect -50 6045 50 6064
rect -50 5026 50 5045
rect -50 5009 -42 5026
rect 42 5009 50 5026
rect -50 5001 50 5009
rect -50 4972 50 4980
rect -50 4955 -42 4972
rect 42 4955 50 4972
rect -50 4936 50 4955
rect -50 3917 50 3936
rect -50 3900 -42 3917
rect 42 3900 50 3917
rect -50 3892 50 3900
rect -50 3863 50 3871
rect -50 3846 -42 3863
rect 42 3846 50 3863
rect -50 3827 50 3846
rect -50 2808 50 2827
rect -50 2791 -42 2808
rect 42 2791 50 2808
rect -50 2783 50 2791
rect -50 2754 50 2762
rect -50 2737 -42 2754
rect 42 2737 50 2754
rect -50 2718 50 2737
rect -50 1699 50 1718
rect -50 1682 -42 1699
rect 42 1682 50 1699
rect -50 1674 50 1682
rect -50 1645 50 1653
rect -50 1628 -42 1645
rect 42 1628 50 1645
rect -50 1609 50 1628
rect -50 590 50 609
rect -50 573 -42 590
rect 42 573 50 590
rect -50 565 50 573
rect -50 536 50 544
rect -50 519 -42 536
rect 42 519 50 536
rect -50 500 50 519
rect -50 -519 50 -500
rect -50 -536 -42 -519
rect 42 -536 50 -519
rect -50 -544 50 -536
rect -50 -573 50 -565
rect -50 -590 -42 -573
rect 42 -590 50 -573
rect -50 -609 50 -590
rect -50 -1628 50 -1609
rect -50 -1645 -42 -1628
rect 42 -1645 50 -1628
rect -50 -1653 50 -1645
rect -50 -1682 50 -1674
rect -50 -1699 -42 -1682
rect 42 -1699 50 -1682
rect -50 -1718 50 -1699
rect -50 -2737 50 -2718
rect -50 -2754 -42 -2737
rect 42 -2754 50 -2737
rect -50 -2762 50 -2754
rect -50 -2791 50 -2783
rect -50 -2808 -42 -2791
rect 42 -2808 50 -2791
rect -50 -2827 50 -2808
rect -50 -3846 50 -3827
rect -50 -3863 -42 -3846
rect 42 -3863 50 -3846
rect -50 -3871 50 -3863
rect -50 -3900 50 -3892
rect -50 -3917 -42 -3900
rect 42 -3917 50 -3900
rect -50 -3936 50 -3917
rect -50 -4955 50 -4936
rect -50 -4972 -42 -4955
rect 42 -4972 50 -4955
rect -50 -4980 50 -4972
rect -50 -5009 50 -5001
rect -50 -5026 -42 -5009
rect 42 -5026 50 -5009
rect -50 -5045 50 -5026
rect -50 -6064 50 -6045
rect -50 -6081 -42 -6064
rect 42 -6081 50 -6064
rect -50 -6089 50 -6081
rect -50 -6118 50 -6110
rect -50 -6135 -42 -6118
rect 42 -6135 50 -6118
rect -50 -6154 50 -6135
rect -50 -7173 50 -7154
rect -50 -7190 -42 -7173
rect 42 -7190 50 -7173
rect -50 -7198 50 -7190
rect -50 -7227 50 -7219
rect -50 -7244 -42 -7227
rect 42 -7244 50 -7227
rect -50 -7263 50 -7244
rect -50 -8282 50 -8263
rect -50 -8299 -42 -8282
rect 42 -8299 50 -8282
rect -50 -8307 50 -8299
<< polycont >>
rect -42 8282 42 8299
rect -42 7227 42 7244
rect -42 7173 42 7190
rect -42 6118 42 6135
rect -42 6064 42 6081
rect -42 5009 42 5026
rect -42 4955 42 4972
rect -42 3900 42 3917
rect -42 3846 42 3863
rect -42 2791 42 2808
rect -42 2737 42 2754
rect -42 1682 42 1699
rect -42 1628 42 1645
rect -42 573 42 590
rect -42 519 42 536
rect -42 -536 42 -519
rect -42 -590 42 -573
rect -42 -1645 42 -1628
rect -42 -1699 42 -1682
rect -42 -2754 42 -2737
rect -42 -2808 42 -2791
rect -42 -3863 42 -3846
rect -42 -3917 42 -3900
rect -42 -4972 42 -4955
rect -42 -5026 42 -5009
rect -42 -6081 42 -6064
rect -42 -6135 42 -6118
rect -42 -7190 42 -7173
rect -42 -7244 42 -7227
rect -42 -8299 42 -8282
<< locali >>
rect -130 8333 -82 8350
rect 82 8333 130 8350
rect -130 8302 -113 8333
rect 113 8302 130 8333
rect -50 8282 -42 8299
rect 42 8282 50 8299
rect -73 8257 -56 8265
rect -73 7261 -56 7269
rect 56 8257 73 8265
rect 56 7261 73 7269
rect -50 7227 -42 7244
rect 42 7227 50 7244
rect -50 7173 -42 7190
rect 42 7173 50 7190
rect -73 7148 -56 7156
rect -73 6152 -56 6160
rect 56 7148 73 7156
rect 56 6152 73 6160
rect -50 6118 -42 6135
rect 42 6118 50 6135
rect -50 6064 -42 6081
rect 42 6064 50 6081
rect -73 6039 -56 6047
rect -73 5043 -56 5051
rect 56 6039 73 6047
rect 56 5043 73 5051
rect -50 5009 -42 5026
rect 42 5009 50 5026
rect -50 4955 -42 4972
rect 42 4955 50 4972
rect -73 4930 -56 4938
rect -73 3934 -56 3942
rect 56 4930 73 4938
rect 56 3934 73 3942
rect -50 3900 -42 3917
rect 42 3900 50 3917
rect -50 3846 -42 3863
rect 42 3846 50 3863
rect -73 3821 -56 3829
rect -73 2825 -56 2833
rect 56 3821 73 3829
rect 56 2825 73 2833
rect -50 2791 -42 2808
rect 42 2791 50 2808
rect -50 2737 -42 2754
rect 42 2737 50 2754
rect -73 2712 -56 2720
rect -73 1716 -56 1724
rect 56 2712 73 2720
rect 56 1716 73 1724
rect -50 1682 -42 1699
rect 42 1682 50 1699
rect -50 1628 -42 1645
rect 42 1628 50 1645
rect -73 1603 -56 1611
rect -73 607 -56 615
rect 56 1603 73 1611
rect 56 607 73 615
rect -50 573 -42 590
rect 42 573 50 590
rect -50 519 -42 536
rect 42 519 50 536
rect -73 494 -56 502
rect -73 -502 -56 -494
rect 56 494 73 502
rect 56 -502 73 -494
rect -50 -536 -42 -519
rect 42 -536 50 -519
rect -50 -590 -42 -573
rect 42 -590 50 -573
rect -73 -615 -56 -607
rect -73 -1611 -56 -1603
rect 56 -615 73 -607
rect 56 -1611 73 -1603
rect -50 -1645 -42 -1628
rect 42 -1645 50 -1628
rect -50 -1699 -42 -1682
rect 42 -1699 50 -1682
rect -73 -1724 -56 -1716
rect -73 -2720 -56 -2712
rect 56 -1724 73 -1716
rect 56 -2720 73 -2712
rect -50 -2754 -42 -2737
rect 42 -2754 50 -2737
rect -50 -2808 -42 -2791
rect 42 -2808 50 -2791
rect -73 -2833 -56 -2825
rect -73 -3829 -56 -3821
rect 56 -2833 73 -2825
rect 56 -3829 73 -3821
rect -50 -3863 -42 -3846
rect 42 -3863 50 -3846
rect -50 -3917 -42 -3900
rect 42 -3917 50 -3900
rect -73 -3942 -56 -3934
rect -73 -4938 -56 -4930
rect 56 -3942 73 -3934
rect 56 -4938 73 -4930
rect -50 -4972 -42 -4955
rect 42 -4972 50 -4955
rect -50 -5026 -42 -5009
rect 42 -5026 50 -5009
rect -73 -5051 -56 -5043
rect -73 -6047 -56 -6039
rect 56 -5051 73 -5043
rect 56 -6047 73 -6039
rect -50 -6081 -42 -6064
rect 42 -6081 50 -6064
rect -50 -6135 -42 -6118
rect 42 -6135 50 -6118
rect -73 -6160 -56 -6152
rect -73 -7156 -56 -7148
rect 56 -6160 73 -6152
rect 56 -7156 73 -7148
rect -50 -7190 -42 -7173
rect 42 -7190 50 -7173
rect -50 -7244 -42 -7227
rect 42 -7244 50 -7227
rect -73 -7269 -56 -7261
rect -73 -8265 -56 -8257
rect 56 -7269 73 -7261
rect 56 -8265 73 -8257
rect -50 -8299 -42 -8282
rect 42 -8299 50 -8282
rect -130 -8333 -113 -8302
rect 113 -8333 130 -8302
rect -130 -8350 -82 -8333
rect 82 -8350 130 -8333
<< viali >>
rect -42 8282 42 8299
rect -73 7269 -56 8257
rect 56 7269 73 8257
rect -42 7227 42 7244
rect -42 7173 42 7190
rect -73 6160 -56 7148
rect 56 6160 73 7148
rect -42 6118 42 6135
rect -42 6064 42 6081
rect -73 5051 -56 6039
rect 56 5051 73 6039
rect -42 5009 42 5026
rect -42 4955 42 4972
rect -73 3942 -56 4930
rect 56 3942 73 4930
rect -42 3900 42 3917
rect -42 3846 42 3863
rect -73 2833 -56 3821
rect 56 2833 73 3821
rect -42 2791 42 2808
rect -42 2737 42 2754
rect -73 1724 -56 2712
rect 56 1724 73 2712
rect -42 1682 42 1699
rect -42 1628 42 1645
rect -73 615 -56 1603
rect 56 615 73 1603
rect -42 573 42 590
rect -42 519 42 536
rect -73 -494 -56 494
rect 56 -494 73 494
rect -42 -536 42 -519
rect -42 -590 42 -573
rect -73 -1603 -56 -615
rect 56 -1603 73 -615
rect -42 -1645 42 -1628
rect -42 -1699 42 -1682
rect -73 -2712 -56 -1724
rect 56 -2712 73 -1724
rect -42 -2754 42 -2737
rect -42 -2808 42 -2791
rect -73 -3821 -56 -2833
rect 56 -3821 73 -2833
rect -42 -3863 42 -3846
rect -42 -3917 42 -3900
rect -73 -4930 -56 -3942
rect 56 -4930 73 -3942
rect -42 -4972 42 -4955
rect -42 -5026 42 -5009
rect -73 -6039 -56 -5051
rect 56 -6039 73 -5051
rect -42 -6081 42 -6064
rect -42 -6135 42 -6118
rect -73 -7148 -56 -6160
rect 56 -7148 73 -6160
rect -42 -7190 42 -7173
rect -42 -7244 42 -7227
rect -73 -8257 -56 -7269
rect 56 -8257 73 -7269
rect -42 -8299 42 -8282
<< metal1 >>
rect -48 8299 48 8302
rect -48 8282 -42 8299
rect 42 8282 48 8299
rect -48 8279 48 8282
rect -76 8257 -53 8263
rect -76 7269 -73 8257
rect -56 7269 -53 8257
rect -76 7263 -53 7269
rect 53 8257 76 8263
rect 53 7269 56 8257
rect 73 7269 76 8257
rect 53 7263 76 7269
rect -48 7244 48 7247
rect -48 7227 -42 7244
rect 42 7227 48 7244
rect -48 7224 48 7227
rect -48 7190 48 7193
rect -48 7173 -42 7190
rect 42 7173 48 7190
rect -48 7170 48 7173
rect -76 7148 -53 7154
rect -76 6160 -73 7148
rect -56 6160 -53 7148
rect -76 6154 -53 6160
rect 53 7148 76 7154
rect 53 6160 56 7148
rect 73 6160 76 7148
rect 53 6154 76 6160
rect -48 6135 48 6138
rect -48 6118 -42 6135
rect 42 6118 48 6135
rect -48 6115 48 6118
rect -48 6081 48 6084
rect -48 6064 -42 6081
rect 42 6064 48 6081
rect -48 6061 48 6064
rect -76 6039 -53 6045
rect -76 5051 -73 6039
rect -56 5051 -53 6039
rect -76 5045 -53 5051
rect 53 6039 76 6045
rect 53 5051 56 6039
rect 73 5051 76 6039
rect 53 5045 76 5051
rect -48 5026 48 5029
rect -48 5009 -42 5026
rect 42 5009 48 5026
rect -48 5006 48 5009
rect -48 4972 48 4975
rect -48 4955 -42 4972
rect 42 4955 48 4972
rect -48 4952 48 4955
rect -76 4930 -53 4936
rect -76 3942 -73 4930
rect -56 3942 -53 4930
rect -76 3936 -53 3942
rect 53 4930 76 4936
rect 53 3942 56 4930
rect 73 3942 76 4930
rect 53 3936 76 3942
rect -48 3917 48 3920
rect -48 3900 -42 3917
rect 42 3900 48 3917
rect -48 3897 48 3900
rect -48 3863 48 3866
rect -48 3846 -42 3863
rect 42 3846 48 3863
rect -48 3843 48 3846
rect -76 3821 -53 3827
rect -76 2833 -73 3821
rect -56 2833 -53 3821
rect -76 2827 -53 2833
rect 53 3821 76 3827
rect 53 2833 56 3821
rect 73 2833 76 3821
rect 53 2827 76 2833
rect -48 2808 48 2811
rect -48 2791 -42 2808
rect 42 2791 48 2808
rect -48 2788 48 2791
rect -48 2754 48 2757
rect -48 2737 -42 2754
rect 42 2737 48 2754
rect -48 2734 48 2737
rect -76 2712 -53 2718
rect -76 1724 -73 2712
rect -56 1724 -53 2712
rect -76 1718 -53 1724
rect 53 2712 76 2718
rect 53 1724 56 2712
rect 73 1724 76 2712
rect 53 1718 76 1724
rect -48 1699 48 1702
rect -48 1682 -42 1699
rect 42 1682 48 1699
rect -48 1679 48 1682
rect -48 1645 48 1648
rect -48 1628 -42 1645
rect 42 1628 48 1645
rect -48 1625 48 1628
rect -76 1603 -53 1609
rect -76 615 -73 1603
rect -56 615 -53 1603
rect -76 609 -53 615
rect 53 1603 76 1609
rect 53 615 56 1603
rect 73 615 76 1603
rect 53 609 76 615
rect -48 590 48 593
rect -48 573 -42 590
rect 42 573 48 590
rect -48 570 48 573
rect -48 536 48 539
rect -48 519 -42 536
rect 42 519 48 536
rect -48 516 48 519
rect -76 494 -53 500
rect -76 -494 -73 494
rect -56 -494 -53 494
rect -76 -500 -53 -494
rect 53 494 76 500
rect 53 -494 56 494
rect 73 -494 76 494
rect 53 -500 76 -494
rect -48 -519 48 -516
rect -48 -536 -42 -519
rect 42 -536 48 -519
rect -48 -539 48 -536
rect -48 -573 48 -570
rect -48 -590 -42 -573
rect 42 -590 48 -573
rect -48 -593 48 -590
rect -76 -615 -53 -609
rect -76 -1603 -73 -615
rect -56 -1603 -53 -615
rect -76 -1609 -53 -1603
rect 53 -615 76 -609
rect 53 -1603 56 -615
rect 73 -1603 76 -615
rect 53 -1609 76 -1603
rect -48 -1628 48 -1625
rect -48 -1645 -42 -1628
rect 42 -1645 48 -1628
rect -48 -1648 48 -1645
rect -48 -1682 48 -1679
rect -48 -1699 -42 -1682
rect 42 -1699 48 -1682
rect -48 -1702 48 -1699
rect -76 -1724 -53 -1718
rect -76 -2712 -73 -1724
rect -56 -2712 -53 -1724
rect -76 -2718 -53 -2712
rect 53 -1724 76 -1718
rect 53 -2712 56 -1724
rect 73 -2712 76 -1724
rect 53 -2718 76 -2712
rect -48 -2737 48 -2734
rect -48 -2754 -42 -2737
rect 42 -2754 48 -2737
rect -48 -2757 48 -2754
rect -48 -2791 48 -2788
rect -48 -2808 -42 -2791
rect 42 -2808 48 -2791
rect -48 -2811 48 -2808
rect -76 -2833 -53 -2827
rect -76 -3821 -73 -2833
rect -56 -3821 -53 -2833
rect -76 -3827 -53 -3821
rect 53 -2833 76 -2827
rect 53 -3821 56 -2833
rect 73 -3821 76 -2833
rect 53 -3827 76 -3821
rect -48 -3846 48 -3843
rect -48 -3863 -42 -3846
rect 42 -3863 48 -3846
rect -48 -3866 48 -3863
rect -48 -3900 48 -3897
rect -48 -3917 -42 -3900
rect 42 -3917 48 -3900
rect -48 -3920 48 -3917
rect -76 -3942 -53 -3936
rect -76 -4930 -73 -3942
rect -56 -4930 -53 -3942
rect -76 -4936 -53 -4930
rect 53 -3942 76 -3936
rect 53 -4930 56 -3942
rect 73 -4930 76 -3942
rect 53 -4936 76 -4930
rect -48 -4955 48 -4952
rect -48 -4972 -42 -4955
rect 42 -4972 48 -4955
rect -48 -4975 48 -4972
rect -48 -5009 48 -5006
rect -48 -5026 -42 -5009
rect 42 -5026 48 -5009
rect -48 -5029 48 -5026
rect -76 -5051 -53 -5045
rect -76 -6039 -73 -5051
rect -56 -6039 -53 -5051
rect -76 -6045 -53 -6039
rect 53 -5051 76 -5045
rect 53 -6039 56 -5051
rect 73 -6039 76 -5051
rect 53 -6045 76 -6039
rect -48 -6064 48 -6061
rect -48 -6081 -42 -6064
rect 42 -6081 48 -6064
rect -48 -6084 48 -6081
rect -48 -6118 48 -6115
rect -48 -6135 -42 -6118
rect 42 -6135 48 -6118
rect -48 -6138 48 -6135
rect -76 -6160 -53 -6154
rect -76 -7148 -73 -6160
rect -56 -7148 -53 -6160
rect -76 -7154 -53 -7148
rect 53 -6160 76 -6154
rect 53 -7148 56 -6160
rect 73 -7148 76 -6160
rect 53 -7154 76 -7148
rect -48 -7173 48 -7170
rect -48 -7190 -42 -7173
rect 42 -7190 48 -7173
rect -48 -7193 48 -7190
rect -48 -7227 48 -7224
rect -48 -7244 -42 -7227
rect 42 -7244 48 -7227
rect -48 -7247 48 -7244
rect -76 -7269 -53 -7263
rect -76 -8257 -73 -7269
rect -56 -8257 -53 -7269
rect -76 -8263 -53 -8257
rect 53 -7269 76 -7263
rect 53 -8257 56 -7269
rect 73 -8257 76 -7269
rect 53 -8263 76 -8257
rect -48 -8282 48 -8279
rect -48 -8299 -42 -8282
rect 42 -8299 48 -8282
rect -48 -8302 48 -8299
<< properties >>
string FIXED_BBOX -121 -8341 121 8341
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 15 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
