** sch_path: /foss/designs/sim/tb_tt06_tempsens.sch
**.subckt tb_tt06_tempsens
VDD1 VDD GND 1.8
VCLK clk GND 0 pulse(0 1.8 0 1n 1n {0.5/fclk} {1/fclk})
VRES rstn GND 1.8 pwl(0 1.8 0.5u 1.8 0.501u 0)
x1 clk VDD rstn VDD VDD VDD VDD VDD GND GND GND GND net4 net3 net1 st11 deb0 deb1 deb2 deb3 st1 st2 st3 st5 st6 st7 daccode st10
+ VDD st8 net5 st0 daccode net7 net2 prechrgn net8 st9 net6 VDD VDD st4 VDD VDD GND tt_um_hpretl_tt06_tempsens
C1 st7 GND 10f m=1
C3 st1 GND 10f m=1
C4 st0 GND 10f m=1
C2 st3 GND 10f m=1
C5 st2 GND 10f m=1
C6 st5 GND 10f m=1
C7 st4 GND 10f m=1
C8 st6 GND 10f m=1
C9 deb3 GND 10f m=1
C10 st9 GND 10f m=1
C11 st8 GND 10f m=1
C12 st11 GND 10f m=1
C13 st10 GND 10f m=1
C14 deb1 GND 10f m=1
C15 deb0 GND 10f m=1
C16 deb2 GND 10f m=1
C17 net1 GND 10f m=1
C18 net7 GND 10f m=1
C19 net8 GND 10f m=1
C20 net5 GND 10f m=1
C21 net6 GND 10f m=1
C22 net3 GND 10f m=1
C23 net4 GND 10f m=1
C24 net2 GND 10f m=1
.save v(deb0)
.save v(rstn)
.save v(clk)
VDAC daccode GND 1.8 pwl(0 1.8 1u 1.8 1.001u 0)
.save v(daccode)
VDAC1 prechrgn GND 1.8 pwl(0 0 1.1u 0 1.101u 1.8)
.save v(prechrgn)
**** begin user architecture code



* ngspice commands
****************

****************
* Misc
****************
.param fclk=10MEG
.options method=gear maxord=2
.temp 30

.save x1.ts.ts_core.dac_vout_ana_
.save x1.ts.ts_core.dcdel_capnode_ana_

.control
set num_threads=6
tran 5u 250u

*exit
.endc




** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  tt_um_hpretl_tt06_tempsens.sym # of pins=45
** sym_path: /foss/designs/sim/tt_um_hpretl_tt06_tempsens.sym
.include tt_um_hpretl_tt06_tempsens.pex.spice
.GLOBAL VDD
.GLOBAL GND
.end
