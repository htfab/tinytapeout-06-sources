module longest_run_of_ones_core (
  clk, rst_n, valid_rsc_dat, valid_triosy_lz, is_random_rsc_dat, is_random_triosy_lz,
      epsilon_rsc_dat, epsilon_triosy_lz
);
  input clk;
  input rst_n;
  output valid_rsc_dat;
  output valid_triosy_lz;
  output is_random_rsc_dat;
  output is_random_triosy_lz;
  input epsilon_rsc_dat;
  output epsilon_triosy_lz;


  // Interconnect Declarations
  reg valid_rsci_idat;
  reg is_random_rsci_idat;
  wire epsilon_rsci_idat;
  wire if_2_if_if_2_if_or_471_tmp;
  wire if_2_aif_2_if_2_aelse_2_and_tmp;
  wire [6:0] mux_7_tmp;
  wire [6:0] mux_6_tmp;
  wire [6:0] mux_5_tmp;
  wire [6:0] mux_4_tmp;
  wire [6:0] mux_1_tmp;
  wire [6:0] acc_tmp;
  wire [7:0] nl_acc_tmp;
  wire and_dcpl;
  wire and_dcpl_3;
  wire and_dcpl_8;
  wire or_dcpl_7;
  wire or_dcpl_10;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_23;
  wire or_dcpl_28;
  wire or_dcpl_31;
  wire and_dcpl_10;
  wire and_dcpl_12;
  wire and_dcpl_13;
  wire and_dcpl_16;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_22;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire or_tmp_3;
  wire mux_tmp;
  wire and_dcpl_28;
  wire or_dcpl_38;
  wire mux_tmp_11;
  wire and_dcpl_30;
  wire mux_tmp_22;
  wire or_tmp_35;
  wire and_dcpl_32;
  wire not_tmp_52;
  wire mux_tmp_34;
  wire and_dcpl_34;
  wire or_tmp_55;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_41;
  wire and_dcpl_42;
  wire and_dcpl_45;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire not_tmp_66;
  wire and_dcpl_55;
  wire and_dcpl_58;
  wire and_dcpl_60;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_69;
  wire or_tmp_75;
  wire mux_tmp_63;
  wire mux_tmp_65;
  wire mux_tmp_66;
  wire and_dcpl_71;
  wire or_tmp_83;
  wire mux_tmp_68;
  wire and_dcpl_73;
  wire mux_tmp_70;
  wire and_dcpl_75;
  wire and_dcpl_77;
  wire and_dcpl_87;
  wire and_dcpl_92;
  wire and_dcpl_96;
  wire and_dcpl_110;
  wire and_dcpl_121;
  wire if_2_oif_13_aelse_2_nor_cse_1;
  wire if_2_oif_13_aelse_1_nor_2;
  wire if_2_oif_468_aelse_nor_2;
  wire if_2_if_2_if_nor_cse_sva_1;
  wire if_2_oif_7_aelse_2_nor_cse_1;
  wire if_2_oif_12_aelse_1_nor_2;
  wire if_2_oif_2_aelse_2_nor_cse_1;
  wire if_2_oif_11_aelse_1_nor_2;
  wire if_2_oif_1_aelse_2_nor_cse_1;
  wire if_2_aelse_1_nor_cse_1;
  wire if_2_oif_aelse_2_nor_cse_1;
  wire if_2_oif_9_aelse_1_nor_2;
  wire if_2_aelse_2_nor_cse_1;
  wire if_2_oif_8_aelse_1_nor_2;
  wire if_2_oif_465_aelse_nor_2;
  wire if_2_aelse_nor_cse_1;
  wire if_1_switch_lp_equal_tmp_2;
  wire if_1_switch_lp_equal_tmp_3;
  reg [6:0] n_sva;
  wire [6:0] nu_3_sva_dfm_1_mx0;
  wire if_2_oif_13_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_13_land_1_lpi_1_dfm;
  wire [3:0] nu_2_sva_dfm_1_mx0_6_3;
  wire nu_1_sva_dfm_1_mx1_2;
  wire [1:0] nu_1_sva_dfm_1_mx0_1_0;
  wire if_2_oif_12_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_12_land_1_lpi_1_dfm;
  wire nu_2_sva_dfm_1_mx1_2;
  wire nu_2_sva_dfm_1_mx0_1;
  wire nu_2_sva_dfm_1_mx1_0;
  wire if_2_oif_11_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_11_land_1_lpi_1_dfm;
  wire if_2_oif_10_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_10_land_1_lpi_1_dfm;
  wire if_2_oif_9_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_9_land_1_lpi_1_dfm;
  wire if_2_oif_8_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_8_land_1_lpi_1_dfm;
  wire if_2_oif_7_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_7_land_1_lpi_1_dfm;
  wire if_2_oif_6_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_6_land_1_lpi_1_dfm;
  wire if_2_oif_5_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_5_land_1_lpi_1_dfm;
  wire if_2_oif_4_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_4_land_1_lpi_1_dfm;
  wire if_2_oif_3_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_3_land_1_lpi_1_dfm;
  wire if_2_oif_2_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_2_land_1_lpi_1_dfm;
  wire if_2_oif_1_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_1_land_1_lpi_1_dfm;
  wire [3:0] nu_1_sva_dfm_1_mx0_6_3;
  wire [6:0] nu_0_sva_dfm_1_mx0;
  wire [6:0] v_n_obs_sva_dfm_1_mx0;
  reg reg_epsilon_triosy_obj_ld_cse;
  wire or_40_cse;
  wire and_134_cse;
  wire nand_22_cse;
  wire or_44_cse;
  wire nor_19_cse;
  wire nand_23_cse;
  wire or_36_cse;
  wire or_81_cse;
  wire or_69_cse;
  wire or_85_cse;
  wire nor_25_cse;
  wire if_2_oif_470_aelse_1_nor_2;
  wire if_2_oelse_447_nor_3;
  wire if_2_oif_20_aelse_2_nor_cse_1;
  wire if_2_oif_472_aelse_1_nor_2;
  wire if_2_oif_45_aelse_nor_2;
  wire if_2_oif_44_aelse_nor_2;
  wire if_2_oif_104_aelse_nor_2;
  wire if_2_oif_21_aelse_nor_2;
  wire if_2_oelse_409_nor_3;
  wire if_2_oif_471_aelse_nor_2;
  wire if_2_oelse_409_if_2_oelse_409_nor_2;
  wire if_2_oif_27_aelse_nor_2;
  wire if_2_oelse_361_nor_3;
  wire if_2_oelse_361_if_2_oelse_361_nor_2;
  wire if_2_oif_33_aelse_nor_2;
  wire if_2_oelse_302_nor_3;
  wire if_2_oelse_302_if_2_oelse_302_nor_2;
  wire if_2_oif_39_aelse_nor_2;
  wire if_2_oelse_239_nor_3;
  wire if_2_oelse_239_if_2_oelse_239_nor_2;
  wire if_2_oelse_173_nor_3;
  wire if_2_oif_49_aelse_2_nor_cse_1;
  wire if_2_oif_43_aelse_nor_2;
  wire if_2_oelse_104_nor_3;
  wire if_2_oif_115_aelse_1_nor_2;
  wire if_2_oelse_44_nor_3;
  wire if_2_oif_14_land_1_lpi_1_dfm_mx0w0;
  reg if_2_oif_14_land_1_lpi_1_dfm;
  reg [6:0] run_sva;
  reg [6:0] v_n_obs_sva;
  reg [6:0] nu_1_sva;
  reg [6:0] nu_2_sva;
  reg [6:0] nu_0_sva;
  reg [6:0] nu_3_sva;
  reg if_2_lor_471_lpi_1_dfm_1;
  reg if_2_oif_472_land_1_lpi_1_dfm;
  wire [6:0] run_sva_2;
  wire [7:0] nl_run_sva_2;
  wire [6:0] asn_25_mx0w1;
  wire [7:0] nl_asn_25_mx0w1;
  wire [6:0] asn_20_mx0w0;
  wire [7:0] nl_asn_20_mx0w0;
  wire [6:0] nu_3_sva_dfm_1_mx1;
  wire if_1_switch_lp_nor_tmp_1;
  wire [6:0] asn_22_mx0w0;
  wire [7:0] nl_asn_22_mx0w0;
  wire [6:0] asn_24_mx0w0;
  wire [7:0] nl_asn_24_mx0w0;
  wire if_2_oif_472_land_1_lpi_1_dfm_mx0;
  wire if_2_lor_471_lpi_1_dfm_1_mx0;
  wire unequal_tmp_2;
  wire unequal_tmp_3;
  wire and_149_cse;
  wire and_178_cse;
  wire if_if_acc_itm_7;

  wire mux_93_nl;
  wire nor_56_nl;
  wire nor_57_nl;
  wire mux_94_nl;
  wire nor_58_nl;
  wire nor_59_nl;
  wire mux_95_nl;
  wire nor_60_nl;
  wire nor_61_nl;
  wire mux_96_nl;
  wire or_1545_nl;
  wire or_1544_nl;
  wire nand_35_nl;
  wire[7:0] if_if_acc_nl;
  wire[8:0] nl_if_if_acc_nl;
  wire and_16_nl;
  wire or_10_nl;
  wire if_2_oif_472_aif_1_if_2_oif_472_aelse_1_and_nl;
  wire or_33_nl;
  wire if_2_oif_14_aelse_1_mux_nl;
  wire if_2_oif_13_aelse_1_mux_nl;
  wire if_2_oif_12_aelse_1_mux_nl;
  wire if_2_oif_11_aelse_1_mux_nl;
  wire if_2_oif_10_aelse_1_mux_nl;
  wire if_2_oif_9_aelse_1_mux_nl;
  wire if_2_oif_8_aelse_1_mux_nl;
  wire if_2_oif_7_aelse_1_mux_nl;
  wire if_2_oif_6_aelse_1_mux_nl;
  wire if_2_oif_5_aelse_1_mux_nl;
  wire if_2_oif_4_aelse_1_mux_nl;
  wire if_2_oif_3_aelse_1_mux_nl;
  wire if_2_oif_2_aelse_1_mux_nl;
  wire if_2_oif_1_aelse_1_mux_nl;
  wire or_35_nl;
  wire and_12_nl;
  wire and_11_nl;
  wire and_10_nl;
  wire or_nl;
  wire mux_24_nl;
  wire and_nl;
  wire mux_23_nl;
  wire nor_18_nl;
  wire mux_22_nl;
  wire mux_21_nl;
  wire and_135_nl;
  wire mux_20_nl;
  wire mux_19_nl;
  wire mux_18_nl;
  wire nor_20_nl;
  wire mux_17_nl;
  wire mux_16_nl;
  wire mux_15_nl;
  wire or_38_nl;
  wire mux_35_nl;
  wire and_137_nl;
  wire mux_34_nl;
  wire nor_21_nl;
  wire mux_33_nl;
  wire mux_32_nl;
  wire and_138_nl;
  wire mux_31_nl;
  wire mux_30_nl;
  wire mux_29_nl;
  wire nor_23_nl;
  wire mux_28_nl;
  wire mux_27_nl;
  wire mux_26_nl;
  wire or_56_nl;
  wire mux_45_nl;
  wire mux_44_nl;
  wire mux_43_nl;
  wire nand_6_nl;
  wire mux_42_nl;
  wire mux_41_nl;
  wire or_79_nl;
  wire mux_40_nl;
  wire mux_39_nl;
  wire mux_38_nl;
  wire mux_37_nl;
  wire or_73_nl;
  wire or_71_nl;
  wire nor_24_nl;
  wire nand_28_nl;
  wire or_89_nl;
  wire mux_53_nl;
  wire mux_52_nl;
  wire mux_51_nl;
  wire mux_50_nl;
  wire nand_8_nl;
  wire mux_49_nl;
  wire mux_47_nl;
  wire nand_7_nl;
  wire mux_62_nl;
  wire nor_27_nl;
  wire mux_61_nl;
  wire mux_60_nl;
  wire mux_59_nl;
  wire and_143_nl;
  wire mux_58_nl;
  wire nand_29_nl;
  wire mux_57_nl;
  wire nand_30_nl;
  wire and_144_nl;
  wire mux_56_nl;
  wire mux_55_nl;
  wire or_101_nl;
  wire or_100_nl;
  wire nor_28_nl;
  wire and_145_nl;
  wire mux_54_nl;
  wire and_142_nl;
  wire nor_26_nl;
  wire mux_69_nl;
  wire mux_68_nl;
  wire mux_67_nl;
  wire mux_66_nl;
  wire or_115_nl;
  wire or_114_nl;
  wire or_113_nl;
  wire mux_65_nl;
  wire mux_63_nl;
  wire or_108_nl;
  wire mux_76_nl;
  wire and_148_nl;
  wire mux_75_nl;
  wire nand_12_nl;
  wire mux_74_nl;
  wire or_125_nl;
  wire mux_73_nl;
  wire mux_72_nl;
  wire mux_71_nl;
  wire or_124_nl;
  wire nor_34_nl;
  wire mux_70_nl;
  wire or_122_nl;
  wire or_120_nl;
  wire nand_34_nl;
  wire or_130_nl;
  wire or_134_nl;
  wire or_133_nl;
  wire mux_81_nl;
  wire mux_78_nl;
  wire mux_83_nl;
  wire mux_85_nl;
  wire mux_86_nl;
  wire or_143_nl;
  wire mux_88_nl;
  wire or_1530_nl;
  wire mux_87_nl;
  wire or_149_nl;
  wire or_147_nl;
  wire or_1531_nl;
  wire mux_89_nl;
  wire or_1532_nl;
  wire or_1533_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_out_v1 #(.rscid(32'sd1),
  .width(32'sd1)) valid_rsci (
      .idat(valid_rsci_idat),
      .dat(valid_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd1)) is_random_rsci (
      .idat(is_random_rsci_idat),
      .dat(is_random_rsc_dat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd1)) epsilon_rsci (
      .dat(epsilon_rsc_dat),
      .idat(epsilon_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) valid_triosy_obj (
      .ld(reg_epsilon_triosy_obj_ld_cse),
      .lz(valid_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) is_random_triosy_obj (
      .ld(reg_epsilon_triosy_obj_ld_cse),
      .lz(is_random_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) epsilon_triosy_obj (
      .ld(reg_epsilon_triosy_obj_ld_cse),
      .lz(epsilon_triosy_lz)
    );
  assign and_149_cse = epsilon_rsci_idat & if_if_acc_itm_7;
  assign and_178_cse = (n_sva[6:3]==4'b1111);
  assign nand_35_nl = ~(epsilon_rsci_idat & if_if_acc_itm_7);
  assign v_n_obs_sva_dfm_1_mx0 = MUX_v_7_2_2(run_sva_2, v_n_obs_sva, nand_35_nl);
  assign nl_run_sva_2 = run_sva + 7'b0000001;
  assign run_sva_2 = nl_run_sva_2[6:0];
  assign nl_if_if_acc_nl = ({1'b1 , v_n_obs_sva}) + conv_u2u_7_8(~ run_sva_2) + 8'b00000001;
  assign if_if_acc_nl = nl_if_if_acc_nl[7:0];
  assign if_if_acc_itm_7 = readslicef_8_1_7(if_if_acc_nl);
  assign nl_asn_25_mx0w1 = nu_0_sva + 7'b0000001;
  assign asn_25_mx0w1 = nl_asn_25_mx0w1[6:0];
  assign and_16_nl = and_dcpl_3 & and_dcpl & (~ (mux_1_tmp[1]));
  assign nu_0_sva_dfm_1_mx0 = MUX_v_7_2_2(nu_0_sva, asn_25_mx0w1, and_16_nl);
  assign nl_asn_20_mx0w0 = nu_3_sva + 7'b0000001;
  assign asn_20_mx0w0 = nl_asn_20_mx0w0[6:0];
  assign nu_3_sva_dfm_1_mx0 = MUX_v_7_2_2(asn_20_mx0w0, nu_3_sva, and_dcpl_8);
  assign or_10_nl = and_dcpl_8 | or_dcpl_7 | (~ (n_sva[0]));
  assign nu_3_sva_dfm_1_mx1 = MUX_v_7_2_2(asn_20_mx0w0, nu_3_sva, or_10_nl);
  assign if_1_switch_lp_nor_tmp_1 = ~((~((v_n_obs_sva_dfm_1_mx0!=7'b0000000))) |
      ((v_n_obs_sva_dfm_1_mx0==7'b0000001)) | if_1_switch_lp_equal_tmp_2 | if_1_switch_lp_equal_tmp_3);
  assign if_1_switch_lp_equal_tmp_2 = (v_n_obs_sva_dfm_1_mx0==7'b0000010);
  assign if_1_switch_lp_equal_tmp_3 = (v_n_obs_sva_dfm_1_mx0==7'b0000011);
  assign nl_asn_22_mx0w0 = nu_2_sva + 7'b0000001;
  assign asn_22_mx0w0 = nl_asn_22_mx0w0[6:0];
  assign nu_2_sva_dfm_1_mx0_6_3 = MUX_v_4_2_2((asn_22_mx0w0[6:3]), (nu_2_sva[6:3]),
      or_dcpl_15);
  assign nu_2_sva_dfm_1_mx0_1 = MUX_s_1_2_2((asn_22_mx0w0[1]), (nu_2_sva[1]), or_dcpl_15);
  assign nu_2_sva_dfm_1_mx1_2 = MUX_s_1_2_2((asn_22_mx0w0[2]), (nu_2_sva[2]), or_dcpl_15);
  assign nu_2_sva_dfm_1_mx1_0 = MUX_s_1_2_2((asn_22_mx0w0[0]), (nu_2_sva[0]), or_dcpl_15);
  assign nl_asn_24_mx0w0 = nu_1_sva + 7'b0000001;
  assign asn_24_mx0w0 = nl_asn_24_mx0w0[6:0];
  assign nu_1_sva_dfm_1_mx0_6_3 = MUX_v_4_2_2((asn_24_mx0w0[6:3]), (nu_1_sva[6:3]),
      or_dcpl_23);
  assign nu_1_sva_dfm_1_mx0_1_0 = MUX_v_2_2_2((asn_24_mx0w0[1:0]), (nu_1_sva[1:0]),
      or_dcpl_23);
  assign nu_1_sva_dfm_1_mx1_2 = MUX_s_1_2_2((asn_24_mx0w0[2]), (nu_1_sva[2]), or_dcpl_23);
  assign if_2_oif_472_aif_1_if_2_oif_472_aelse_1_and_nl = nu_2_sva_dfm_1_mx1_0 &
      if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3;
  assign or_33_nl = or_dcpl_31 | or_dcpl_28 | (~ (n_sva[6])) | if_2_if_if_2_if_or_471_tmp;
  assign if_2_oif_472_land_1_lpi_1_dfm_mx0 = MUX_s_1_2_2(if_2_oif_472_aif_1_if_2_oif_472_aelse_1_and_nl,
      if_2_oif_472_land_1_lpi_1_dfm, or_33_nl);
  assign if_2_oif_14_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_14_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_14_land_1_lpi_1_dfm, and_dcpl_28);
  assign if_2_oif_13_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_13_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_13_land_1_lpi_1_dfm, and_dcpl_30);
  assign if_2_oif_12_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_12_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_12_land_1_lpi_1_dfm, and_dcpl_32);
  assign if_2_oif_11_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_11_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_11_land_1_lpi_1_dfm, and_dcpl_34);
  assign if_2_oif_10_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_10_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_10_land_1_lpi_1_dfm, and_dcpl_36);
  assign if_2_oif_9_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_9_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_9_land_1_lpi_1_dfm, and_dcpl_38);
  assign if_2_oif_8_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_8_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_8_land_1_lpi_1_dfm, and_dcpl_55);
  assign if_2_oif_7_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_7_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_7_land_1_lpi_1_dfm, and_dcpl_71);
  assign if_2_oif_6_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_6_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_6_land_1_lpi_1_dfm, and_dcpl_73);
  assign if_2_oif_5_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_5_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_5_land_1_lpi_1_dfm, and_dcpl_75);
  assign if_2_oif_4_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_4_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_4_land_1_lpi_1_dfm, and_dcpl_77);
  assign if_2_oif_3_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_3_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_3_land_1_lpi_1_dfm, and_dcpl_92);
  assign if_2_oif_2_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_2_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_2_land_1_lpi_1_dfm, and_dcpl_110);
  assign if_2_oif_1_aelse_1_mux_nl = MUX_s_1_2_2(if_2_oif_1_land_1_lpi_1_dfm_mx0w0,
      if_2_oif_1_land_1_lpi_1_dfm, and_dcpl_121);
  assign if_2_if_if_2_if_or_471_tmp = ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3])
      & if_2_oelse_447_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 &
      (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 &
      (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3])
      & if_2_oelse_447_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3])
      & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3])
      & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[3]) & if_2_oelse_447_nor_3) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:0]==3'b111) & if_2_oelse_409_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & if_2_oelse_409_if_2_oelse_409_nor_2)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & if_2_oelse_409_if_2_oelse_409_nor_2)
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 &
      (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oelse_361_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & if_2_oelse_361_if_2_oelse_361_nor_2)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & if_2_oelse_361_if_2_oelse_361_nor_2)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & if_2_oelse_361_if_2_oelse_361_nor_2) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2
      & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) &
      if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~((nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & if_2_oelse_302_if_2_oelse_302_nor_2)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      if_2_oelse_302_if_2_oelse_302_nor_2) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) &
      if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 &
      if_2_aelse_1_nor_cse_1 & if_2_oelse_302_if_2_oelse_302_nor_2) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~((nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[2]) & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & if_2_oelse_239_if_2_oelse_239_nor_2)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & if_2_oelse_239_if_2_oelse_239_nor_2)
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~((nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2
      & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[3])
      & if_2_oif_49_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[3]) & if_2_oif_49_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[3])
      & if_2_oif_49_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oelse_173_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oelse_173_nor_3)
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & nu_1_sva_dfm_1_mx1_2 & if_2_oif_43_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & nu_1_sva_dfm_1_mx1_2 & if_2_oif_43_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & nu_1_sva_dfm_1_mx1_2 & if_2_oif_43_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000)
      | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~(nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~((nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[3])
      & if_2_oif_49_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_115_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[3])
      & if_2_oif_49_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0])
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_115_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_13_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[3])
      & if_2_oif_49_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1]) & if_2_oelse_104_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_104_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[1])
      & if_2_oelse_104_nor_3) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & nu_1_sva_dfm_1_mx1_2 & if_2_oif_43_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & nu_1_sva_dfm_1_mx1_2 & if_2_oif_43_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_39_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)))))
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & (~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_2_sva_dfm_1_mx1_2 | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0 | (~((nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3))))) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3)))) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~((nu_2_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_13_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3))))
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 &
      nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[3]) & if_2_oif_49_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2
      & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[3])
      & if_2_oif_49_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 &
      (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) &
      if_2_oif_2_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_45_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_44_nor_3)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_44_aelse_nor_2 & (nu_0_sva_dfm_1_mx0[0])
      & if_2_oelse_44_nor_3) | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & nu_1_sva_dfm_1_mx1_2 & if_2_oif_43_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_39_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_39_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_39_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | (~((nu_3_sva_dfm_1_mx0!=7'b0000000) | (~(nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)))) | ((nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_33_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 &
      (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_33_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_470_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_27_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_472_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_27_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[1]) & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_8_aelse_1_nor_2 & (nu_1_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_21_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & (nu_1_sva_dfm_1_mx0_6_3[0]) & if_2_oif_21_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[0]) & if_2_oif_20_aelse_2_nor_cse_1 & (nu_2_sva_dfm_1_mx0_6_3[0])
      & if_2_oif_13_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx0_1 & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2
      & if_2_oif_9_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11)
      & if_2_oif_471_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_aelse_2_nor_cse_1 & if_2_oif_14_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[1])
      & if_2_oif_13_aelse_2_nor_cse_1 & if_2_oif_13_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11)
      & if_2_oif_7_aelse_2_nor_cse_1 & if_2_oif_12_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2])
      & if_2_oif_2_aelse_2_nor_cse_1 & if_2_oif_11_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2])
      & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1 & if_2_oif_10_aelse_1_mux_nl)
      | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1 & if_2_oif_9_aelse_1_mux_nl)
      | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1 & if_2_oif_8_aelse_1_mux_nl)
      | ((nu_3_sva_dfm_1_mx0[1:0]==2'b11) & if_2_oif_7_aelse_2_nor_cse_1 & if_2_oif_7_aelse_1_mux_nl)
      | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1 & if_2_oif_6_aelse_1_mux_nl)
      | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0]) & if_2_oif_1_aelse_2_nor_cse_1
      & if_2_oif_5_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11) & if_2_oif_aelse_2_nor_cse_1
      & if_2_oif_4_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & if_2_oif_3_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2]) & if_2_oif_2_aelse_2_nor_cse_1
      & if_2_oif_2_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2]) & (nu_3_sva_dfm_1_mx0[0])
      & if_2_oif_1_aelse_2_nor_cse_1 & if_2_oif_1_aelse_1_mux_nl) | ((nu_3_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oif_aelse_2_nor_cse_1 & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 &
      if_2_if_2_if_nor_cse_sva_1) | if_2_aif_2_if_2_aelse_2_and_tmp;
  assign or_35_nl = or_dcpl_31 | or_dcpl_28 | (~ (n_sva[6]));
  assign if_2_lor_471_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(if_2_if_if_2_if_or_471_tmp, if_2_lor_471_lpi_1_dfm_1,
      or_35_nl);
  assign if_2_oif_14_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx0_1 & if_2_oif_470_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0==2'b11) & if_2_oif_471_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_if_2_if_nor_cse_sva_1 = ~((nu_0_sva_dfm_1_mx0!=7'b0000000));
  assign if_2_oif_13_land_1_lpi_1_dfm_mx0w0 = (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_12_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_11_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_10_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_aelse_1_nor_cse_1 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx0_1);
  assign if_2_oif_9_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1]) & if_2_oif_468_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_8_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx0_1 & nu_2_sva_dfm_1_mx1_0
      & if_2_oif_8_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[1])
      & if_2_oif_468_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_7_land_1_lpi_1_dfm_mx0w0 = (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_6_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_5_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & if_2_oif_11_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_4_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0
      & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0])
      & if_2_oif_465_aelse_nor_2 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_3_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & if_2_oif_9_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & (nu_1_sva_dfm_1_mx0_1_0[0]) & if_2_oif_465_aelse_nor_2
      & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_2_land_1_lpi_1_dfm_mx0w0 = (nu_2_sva_dfm_1_mx0_6_3[0]) & if_2_oif_13_aelse_1_nor_2
      & nu_1_sva_dfm_1_mx1_2 & if_2_aelse_nor_cse_1 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_aelse_nor_cse_1 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000) | (nu_1_sva_dfm_1_mx0_1_0!=2'b00));
  assign if_2_oif_1_land_1_lpi_1_dfm_mx0w0 = nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx0_1
      & nu_2_sva_dfm_1_mx1_0 & if_2_oif_12_aelse_1_nor_2 & nu_1_sva_dfm_1_mx1_2 &
      if_2_aelse_nor_cse_1 & if_2_if_2_if_nor_cse_sva_1;
  assign if_2_oif_20_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6:1]!=6'b000000));
  assign if_2_oif_13_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6]) | (nu_3_sva_dfm_1_mx0[5])
      | (nu_3_sva_dfm_1_mx0[4]) | (nu_3_sva_dfm_1_mx0[3]) | (nu_3_sva_dfm_1_mx0[2])
      | (nu_3_sva_dfm_1_mx0[0]));
  assign if_2_oif_7_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6:2]!=5'b00000));
  assign if_2_oif_2_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6]) | (nu_3_sva_dfm_1_mx0[5])
      | (nu_3_sva_dfm_1_mx0[4]) | (nu_3_sva_dfm_1_mx0[3]) | (nu_3_sva_dfm_1_mx0[1])
      | (nu_3_sva_dfm_1_mx0[0]));
  assign if_2_oif_1_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6]) | (nu_3_sva_dfm_1_mx0[5])
      | (nu_3_sva_dfm_1_mx0[4]) | (nu_3_sva_dfm_1_mx0[3]) | (nu_3_sva_dfm_1_mx0[1]));
  assign if_2_oif_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6]) | (nu_3_sva_dfm_1_mx0[5])
      | (nu_3_sva_dfm_1_mx0[4]) | (nu_3_sva_dfm_1_mx0[3]) | (nu_3_sva_dfm_1_mx0[0]));
  assign if_2_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6:3]!=4'b0000));
  assign if_2_oif_49_aelse_2_nor_cse_1 = ~((nu_3_sva_dfm_1_mx0[6]) | (nu_3_sva_dfm_1_mx0[5])
      | (nu_3_sva_dfm_1_mx0[4]) | (nu_3_sva_dfm_1_mx0[2]) | (nu_3_sva_dfm_1_mx0[1])
      | (nu_3_sva_dfm_1_mx0[0]));
  assign if_2_aif_2_if_2_aelse_2_and_tmp = (nu_3_sva_dfm_1_mx0[2:0]==3'b111) & if_2_aelse_2_nor_cse_1
      & nu_2_sva_dfm_1_mx1_2 & nu_2_sva_dfm_1_mx1_0 & if_2_aelse_1_nor_cse_1 & nu_1_sva_dfm_1_mx1_2
      & if_2_aelse_nor_cse_1 & if_2_if_2_if_nor_cse_sva_1;
  assign unequal_tmp_2 = ~((n_sva==7'b1111111));
  assign nl_acc_tmp = n_sva + 7'b0000001;
  assign acc_tmp = nl_acc_tmp[6:0];
  assign unequal_tmp_3 = ~((n_sva[2:0]==3'b111));
  assign if_2_oelse_44_nor_3 = ~((nu_0_sva_dfm_1_mx0[6:1]!=6'b000000));
  assign if_2_oelse_104_nor_3 = ~((nu_0_sva_dfm_1_mx0[6]) | (nu_0_sva_dfm_1_mx0[5])
      | (nu_0_sva_dfm_1_mx0[4]) | (nu_0_sva_dfm_1_mx0[3]) | (nu_0_sva_dfm_1_mx0[2])
      | (nu_0_sva_dfm_1_mx0[0]));
  assign if_2_oelse_173_nor_3 = ~((nu_0_sva_dfm_1_mx0[6:2]!=5'b00000));
  assign if_2_oelse_239_nor_3 = ~((nu_0_sva_dfm_1_mx0[6]) | (nu_0_sva_dfm_1_mx0[5])
      | (nu_0_sva_dfm_1_mx0[4]) | (nu_0_sva_dfm_1_mx0[3]) | (nu_0_sva_dfm_1_mx0[1])
      | (nu_0_sva_dfm_1_mx0[0]));
  assign if_2_oelse_302_nor_3 = ~((nu_0_sva_dfm_1_mx0[6]) | (nu_0_sva_dfm_1_mx0[5])
      | (nu_0_sva_dfm_1_mx0[4]) | (nu_0_sva_dfm_1_mx0[3]) | (nu_0_sva_dfm_1_mx0[1]));
  assign if_2_oelse_361_nor_3 = ~((nu_0_sva_dfm_1_mx0[6]) | (nu_0_sva_dfm_1_mx0[5])
      | (nu_0_sva_dfm_1_mx0[4]) | (nu_0_sva_dfm_1_mx0[3]) | (nu_0_sva_dfm_1_mx0[0]));
  assign if_2_oelse_409_nor_3 = ~((nu_0_sva_dfm_1_mx0[6:3]!=4'b0000));
  assign if_2_oelse_447_nor_3 = ~((nu_0_sva_dfm_1_mx0[6]) | (nu_0_sva_dfm_1_mx0[5])
      | (nu_0_sva_dfm_1_mx0[4]) | (nu_0_sva_dfm_1_mx0[2]) | (nu_0_sva_dfm_1_mx0[1])
      | (nu_0_sva_dfm_1_mx0[0]));
  assign if_2_oif_468_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000) | (nu_1_sva_dfm_1_mx0_1_0[0]));
  assign if_2_oif_465_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000) | (nu_1_sva_dfm_1_mx0_1_0[1]));
  assign if_2_oif_471_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000));
  assign if_2_oif_21_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | nu_1_sva_dfm_1_mx1_2
      | (nu_1_sva_dfm_1_mx0_1_0!=2'b00));
  assign if_2_oif_27_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | nu_1_sva_dfm_1_mx1_2
      | (nu_1_sva_dfm_1_mx0_1_0[1]));
  assign if_2_oif_33_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | nu_1_sva_dfm_1_mx1_2
      | (nu_1_sva_dfm_1_mx0_1_0[0]));
  assign if_2_oif_39_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | nu_1_sva_dfm_1_mx1_2);
  assign if_2_oif_45_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000) | nu_1_sva_dfm_1_mx1_2);
  assign if_2_oif_43_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | (nu_1_sva_dfm_1_mx0_1_0!=2'b00));
  assign if_2_oif_44_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000) | nu_1_sva_dfm_1_mx1_2
      | (nu_1_sva_dfm_1_mx0_1_0[0]));
  assign if_2_oif_104_aelse_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000) | nu_1_sva_dfm_1_mx1_2
      | (nu_1_sva_dfm_1_mx0_1_0[1]));
  assign if_2_oelse_239_if_2_oelse_239_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_1_sva_dfm_1_mx1_2 | (nu_1_sva_dfm_1_mx0_1_0!=2'b00) | (~((nu_0_sva_dfm_1_mx0[2])
      & if_2_oelse_239_nor_3)));
  assign if_2_oelse_302_if_2_oelse_302_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_1_sva_dfm_1_mx1_2 | (nu_1_sva_dfm_1_mx0_1_0!=2'b00) | (~((nu_0_sva_dfm_1_mx0[2])
      & (nu_0_sva_dfm_1_mx0[0]) & if_2_oelse_302_nor_3)));
  assign if_2_oelse_361_if_2_oelse_361_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_1_sva_dfm_1_mx1_2 | (nu_1_sva_dfm_1_mx0_1_0!=2'b00) | (~((nu_0_sva_dfm_1_mx0[2:1]==2'b11)
      & if_2_oelse_361_nor_3)));
  assign if_2_oelse_409_if_2_oelse_409_nor_2 = ~((nu_1_sva_dfm_1_mx0_6_3!=4'b0000)
      | nu_1_sva_dfm_1_mx1_2 | (nu_1_sva_dfm_1_mx0_1_0!=2'b00) | (~((nu_0_sva_dfm_1_mx0[2:0]==3'b111)
      & if_2_oelse_409_nor_3)));
  assign if_2_oif_13_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1 | nu_2_sva_dfm_1_mx1_0);
  assign if_2_oif_12_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000));
  assign if_2_oif_11_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_0);
  assign if_2_oif_9_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx0_1
      | nu_2_sva_dfm_1_mx1_0);
  assign if_2_oif_470_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx1_0);
  assign if_2_oif_8_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2);
  assign if_2_oif_472_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3!=4'b0000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1);
  assign if_2_oif_115_aelse_1_nor_2 = ~((nu_2_sva_dfm_1_mx0_6_3[3:1]!=3'b000) | nu_2_sva_dfm_1_mx1_2
      | nu_2_sva_dfm_1_mx0_1);
  assign and_12_nl = if_1_switch_lp_nor_tmp_1 & (~ unequal_tmp_3);
  assign mux_7_tmp = MUX_v_7_2_2(nu_3_sva, asn_20_mx0w0, and_12_nl);
  assign and_11_nl = if_1_switch_lp_equal_tmp_3 & (~ unequal_tmp_3);
  assign mux_6_tmp = MUX_v_7_2_2(nu_2_sva, asn_22_mx0w0, and_11_nl);
  assign and_10_nl = if_1_switch_lp_equal_tmp_2 & (~ unequal_tmp_3);
  assign mux_5_tmp = MUX_v_7_2_2(nu_1_sva, asn_24_mx0w0, and_10_nl);
  assign or_nl = if_1_switch_lp_equal_tmp_2 | if_1_switch_lp_equal_tmp_3 | if_1_switch_lp_nor_tmp_1
      | unequal_tmp_3;
  assign mux_4_tmp = MUX_v_7_2_2(asn_25_mx0w1, nu_0_sva, or_nl);
  assign mux_1_tmp = MUX_v_7_2_2(v_n_obs_sva, run_sva_2, and_149_cse);
  assign and_dcpl = ~((mux_1_tmp[6:5]!=2'b00));
  assign and_dcpl_3 = ~((mux_1_tmp[4:2]!=3'b000));
  assign and_dcpl_8 = and_dcpl_3 & and_dcpl;
  assign or_dcpl_7 = ~((n_sva[2:1]==2'b11));
  assign or_dcpl_10 = (mux_1_tmp[6]) | (~ (mux_1_tmp[1]));
  assign or_dcpl_14 = (mux_1_tmp[5:2]!=4'b0000);
  assign or_dcpl_15 = or_dcpl_14 | or_dcpl_10 | (~ (mux_1_tmp[0]));
  assign or_dcpl_23 = or_dcpl_14 | or_dcpl_10 | (mux_1_tmp[0]);
  assign or_dcpl_28 = ~((n_sva[5:4]==2'b11));
  assign or_dcpl_31 = or_dcpl_7 | (~((n_sva[0]) & (n_sva[3])));
  assign and_dcpl_10 = ~((mux_7_tmp[5:4]!=2'b00));
  assign and_dcpl_12 = ~((mux_6_tmp[6]) | (mux_7_tmp[3]));
  assign and_dcpl_13 = ~((mux_6_tmp[5:4]!=2'b00));
  assign and_dcpl_16 = ~((mux_5_tmp[5:4]!=2'b00));
  assign and_dcpl_18 = (mux_5_tmp[3:2]==2'b01);
  assign and_dcpl_19 = ~((mux_4_tmp[6:5]!=2'b00));
  assign and_dcpl_22 = and_dcpl_19 & and_dcpl_18 & and_dcpl_16 & (~ (mux_5_tmp[6]))
      & and_dcpl_13 & and_dcpl_12 & and_dcpl_10 & (~ (mux_7_tmp[6]));
  assign and_dcpl_23 = ~((mux_4_tmp[4:3]!=2'b00));
  assign and_dcpl_24 = ~((mux_4_tmp[1:0]!=2'b00));
  assign and_dcpl_25 = and_dcpl_24 & (~ (mux_4_tmp[2]));
  assign and_dcpl_26 = and_dcpl_25 & and_dcpl_23;
  assign or_tmp_3 = (mux_5_tmp[1:0]!=2'b01);
  assign or_40_cse = (mux_5_tmp[1:0]!=2'b10);
  assign mux_tmp = MUX_s_1_2_2(or_40_cse, or_tmp_3, mux_7_tmp[0]);
  assign and_134_cse = (mux_6_tmp[2:0]==3'b111) & (mux_7_tmp[0]) & (mux_5_tmp[1:0]==2'b10);
  assign nand_22_cse = ~((mux_6_tmp[0]) & (mux_7_tmp[0]) & (mux_5_tmp[1:0]==2'b10));
  assign or_44_cse = (mux_5_tmp[1:0]!=2'b00);
  assign nor_19_cse = ~((mux_6_tmp[2:0]!=3'b000) | (mux_7_tmp[0]) | (mux_5_tmp[1:0]!=2'b00));
  assign nand_23_cse = ~((mux_6_tmp[1:0]==2'b11) & (mux_7_tmp[0]) & (mux_5_tmp[1:0]==2'b10));
  assign or_36_cse = (mux_6_tmp[0]) | (mux_7_tmp[0]) | (mux_5_tmp[1:0]!=2'b00);
  assign nor_18_nl = ~((mux_6_tmp[2:0]!=3'b000) | mux_tmp);
  assign mux_23_nl = MUX_s_1_2_2(and_134_cse, nor_18_nl, mux_6_tmp[3]);
  assign and_nl = (mux_7_tmp[1]) & mux_23_nl;
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_3, or_44_cse, mux_7_tmp[0]);
  assign mux_19_nl = MUX_s_1_2_2(mux_tmp, mux_18_nl, mux_6_tmp[0]);
  assign mux_20_nl = MUX_s_1_2_2(nand_22_cse, mux_19_nl, mux_6_tmp[1]);
  assign and_135_nl = (mux_6_tmp[2]) & (~ mux_20_nl);
  assign mux_21_nl = MUX_s_1_2_2(and_135_nl, nor_19_cse, mux_6_tmp[3]);
  assign or_38_nl = (mux_7_tmp[0]) | (mux_5_tmp[1:0]!=2'b01);
  assign mux_15_nl = MUX_s_1_2_2(mux_tmp, or_38_nl, mux_6_tmp[0]);
  assign mux_16_nl = MUX_s_1_2_2(mux_15_nl, or_36_cse, mux_6_tmp[1]);
  assign mux_17_nl = MUX_s_1_2_2(nand_23_cse, mux_16_nl, mux_6_tmp[2]);
  assign nor_20_nl = ~((mux_6_tmp[3]) | mux_17_nl);
  assign mux_22_nl = MUX_s_1_2_2(mux_21_nl, nor_20_nl, mux_7_tmp[1]);
  assign mux_24_nl = MUX_s_1_2_2(and_nl, mux_22_nl, mux_7_tmp[2]);
  assign and_dcpl_28 = mux_24_nl & and_dcpl_26 & and_dcpl_22;
  assign or_dcpl_38 = or_dcpl_31 | or_dcpl_28 | (~ (n_sva[6])) | if_2_aif_2_if_2_aelse_2_and_tmp;
  assign mux_tmp_11 = MUX_s_1_2_2(or_40_cse, or_tmp_3, mux_6_tmp[0]);
  assign nor_21_nl = ~((mux_6_tmp[2:1]!=2'b00) | (~ (mux_7_tmp[0])) | (mux_6_tmp[0])
      | (mux_5_tmp[1:0]!=2'b01));
  assign mux_34_nl = MUX_s_1_2_2(and_134_cse, nor_21_nl, mux_6_tmp[3]);
  assign and_137_nl = (mux_7_tmp[1]) & mux_34_nl;
  assign mux_29_nl = MUX_s_1_2_2(or_tmp_3, or_44_cse, mux_6_tmp[0]);
  assign mux_30_nl = MUX_s_1_2_2(mux_tmp_11, mux_29_nl, mux_7_tmp[0]);
  assign mux_31_nl = MUX_s_1_2_2(nand_22_cse, mux_30_nl, mux_6_tmp[1]);
  assign and_138_nl = (mux_6_tmp[2]) & (~ mux_31_nl);
  assign mux_32_nl = MUX_s_1_2_2(and_138_nl, nor_19_cse, mux_6_tmp[3]);
  assign or_56_nl = (mux_6_tmp[0]) | (mux_5_tmp[1:0]!=2'b01);
  assign mux_26_nl = MUX_s_1_2_2(mux_tmp_11, or_56_nl, mux_7_tmp[0]);
  assign mux_27_nl = MUX_s_1_2_2(mux_26_nl, or_36_cse, mux_6_tmp[1]);
  assign mux_28_nl = MUX_s_1_2_2(nand_23_cse, mux_27_nl, mux_6_tmp[2]);
  assign nor_23_nl = ~((mux_6_tmp[3]) | mux_28_nl);
  assign mux_33_nl = MUX_s_1_2_2(mux_32_nl, nor_23_nl, mux_7_tmp[1]);
  assign mux_35_nl = MUX_s_1_2_2(and_137_nl, mux_33_nl, mux_7_tmp[2]);
  assign and_dcpl_30 = mux_35_nl & and_dcpl_26 & and_dcpl_22;
  assign mux_tmp_22 = MUX_s_1_2_2(or_40_cse, or_44_cse, mux_6_tmp[1]);
  assign or_tmp_35 = (~ (mux_6_tmp[1])) | (mux_5_tmp[1:0]!=2'b01);
  assign or_81_cse = (~ (mux_6_tmp[3])) | (~ (mux_7_tmp[1])) | (mux_6_tmp[2]) | (~
      (mux_7_tmp[0])) | (mux_6_tmp[1:0]!=2'b00) | (mux_5_tmp[1:0]!=2'b01);
  assign or_69_cse = (mux_7_tmp[1]) | (mux_6_tmp[2]) | (mux_7_tmp[0]) | (mux_6_tmp[1:0]!=2'b00)
      | (mux_5_tmp[1:0]!=2'b00);
  assign or_79_nl = (~ (mux_6_tmp[1])) | (mux_5_tmp[1:0]!=2'b10);
  assign mux_41_nl = MUX_s_1_2_2(or_79_nl, or_tmp_35, mux_6_tmp[0]);
  assign mux_40_nl = MUX_s_1_2_2(or_tmp_35, mux_tmp_22, mux_6_tmp[0]);
  assign mux_42_nl = MUX_s_1_2_2(mux_41_nl, mux_40_nl, mux_7_tmp[0]);
  assign nand_6_nl = ~((mux_6_tmp[2]) & (~ mux_42_nl));
  assign or_73_nl = (mux_6_tmp[1]) | (mux_5_tmp[1:0]!=2'b01);
  assign mux_37_nl = MUX_s_1_2_2(mux_tmp_22, or_73_nl, mux_6_tmp[0]);
  assign or_71_nl = (mux_6_tmp[1:0]!=2'b00) | (mux_5_tmp[1:0]!=2'b01);
  assign mux_38_nl = MUX_s_1_2_2(mux_37_nl, or_71_nl, mux_7_tmp[0]);
  assign mux_39_nl = MUX_s_1_2_2(nand_23_cse, mux_38_nl, mux_6_tmp[2]);
  assign mux_43_nl = MUX_s_1_2_2(nand_6_nl, mux_39_nl, mux_7_tmp[1]);
  assign mux_44_nl = MUX_s_1_2_2(mux_43_nl, or_69_cse, mux_6_tmp[3]);
  assign mux_45_nl = MUX_s_1_2_2(or_81_cse, mux_44_nl, mux_7_tmp[2]);
  assign and_dcpl_32 = (~ mux_45_nl) & and_dcpl_26 & and_dcpl_22;
  assign nor_25_cse = ~((mux_5_tmp[1:0]!=2'b00));
  assign nor_24_nl = ~((mux_5_tmp[1:0]!=2'b10));
  assign not_tmp_52 = MUX_s_1_2_2(nor_24_nl, nor_25_cse, mux_6_tmp[1]);
  assign nand_28_nl = ~((mux_6_tmp[2:1]==2'b11) & (mux_5_tmp[1:0]==2'b01));
  assign or_89_nl = (mux_6_tmp[2:1]!=2'b10) | (mux_5_tmp[1:0]!=2'b01);
  assign mux_tmp_34 = MUX_s_1_2_2(nand_28_nl, or_89_nl, mux_7_tmp[1]);
  assign or_85_cse = (mux_6_tmp[2:1]!=2'b01) | (mux_5_tmp[1:0]!=2'b10);
  assign nand_8_nl = ~((mux_7_tmp[1]) & (mux_6_tmp[2]) & not_tmp_52);
  assign mux_50_nl = MUX_s_1_2_2(nand_8_nl, mux_tmp_34, mux_7_tmp[0]);
  assign nand_7_nl = ~((mux_6_tmp[2]) & not_tmp_52);
  assign mux_47_nl = MUX_s_1_2_2(nand_7_nl, or_85_cse, mux_7_tmp[1]);
  assign mux_49_nl = MUX_s_1_2_2(mux_tmp_34, mux_47_nl, mux_7_tmp[0]);
  assign mux_51_nl = MUX_s_1_2_2(mux_50_nl, mux_49_nl, mux_6_tmp[0]);
  assign mux_52_nl = MUX_s_1_2_2(mux_51_nl, or_69_cse, mux_6_tmp[3]);
  assign mux_53_nl = MUX_s_1_2_2(or_81_cse, mux_52_nl, mux_7_tmp[2]);
  assign and_dcpl_34 = (~ mux_53_nl) & and_dcpl_26 & and_dcpl_22;
  assign or_tmp_55 = (~ (mux_6_tmp[1])) | (mux_5_tmp[0]);
  assign nor_27_nl = ~((mux_5_tmp[1]) | (~ (mux_6_tmp[3])) | (~ (mux_7_tmp[1])) |
      (mux_6_tmp[2]) | (~ (mux_7_tmp[0])) | (mux_6_tmp[1:0]!=2'b00) | (~ (mux_5_tmp[0])));
  assign nand_29_nl = ~((mux_6_tmp[1:0]==2'b11) & (mux_5_tmp[0]));
  assign nand_30_nl = ~((mux_6_tmp[1]) & (mux_5_tmp[0]));
  assign mux_57_nl = MUX_s_1_2_2(nand_30_nl, or_tmp_55, mux_6_tmp[0]);
  assign mux_58_nl = MUX_s_1_2_2(nand_29_nl, mux_57_nl, mux_7_tmp[0]);
  assign and_143_nl = (mux_6_tmp[2]) & (~ mux_58_nl);
  assign or_101_nl = (mux_6_tmp[1]) | (~ (mux_5_tmp[0]));
  assign mux_55_nl = MUX_s_1_2_2(or_tmp_55, or_101_nl, mux_6_tmp[0]);
  assign or_100_nl = (mux_6_tmp[1:0]!=2'b00) | (~ (mux_5_tmp[0]));
  assign mux_56_nl = MUX_s_1_2_2(mux_55_nl, or_100_nl, mux_7_tmp[0]);
  assign and_144_nl = (mux_6_tmp[2]) & (~ mux_56_nl);
  assign mux_59_nl = MUX_s_1_2_2(and_143_nl, and_144_nl, mux_7_tmp[1]);
  assign nor_28_nl = ~((mux_7_tmp[1]) | (mux_6_tmp[2]) | (mux_7_tmp[0]) | (mux_6_tmp[1:0]!=2'b00)
      | (mux_5_tmp[0]));
  assign mux_60_nl = MUX_s_1_2_2(mux_59_nl, nor_28_nl, mux_6_tmp[3]);
  assign and_142_nl = (mux_7_tmp[0]) & (mux_6_tmp[1:0]==2'b11) & (~ (mux_5_tmp[0]));
  assign nor_26_nl = ~((mux_7_tmp[0]) | (mux_6_tmp[1:0]!=2'b00) | (mux_5_tmp[0]));
  assign mux_54_nl = MUX_s_1_2_2(and_142_nl, nor_26_nl, mux_6_tmp[2]);
  assign and_145_nl = (~((mux_6_tmp[3]) | (~ (mux_7_tmp[1])))) & mux_54_nl;
  assign mux_61_nl = MUX_s_1_2_2(mux_60_nl, and_145_nl, mux_5_tmp[1]);
  assign mux_62_nl = MUX_s_1_2_2(nor_27_nl, mux_61_nl, mux_7_tmp[2]);
  assign and_dcpl_36 = mux_62_nl & and_dcpl_26 & and_dcpl_22;
  assign or_115_nl = (~ (mux_7_tmp[1])) | (mux_6_tmp[2:1]!=2'b11) | (mux_5_tmp[1:0]!=2'b00);
  assign mux_66_nl = MUX_s_1_2_2(or_115_nl, mux_tmp_34, mux_7_tmp[0]);
  assign or_114_nl = (mux_7_tmp[1:0]!=2'b00) | (mux_6_tmp[2:1]!=2'b00) | (mux_5_tmp[1:0]!=2'b00);
  assign mux_67_nl = MUX_s_1_2_2(mux_66_nl, or_114_nl, mux_6_tmp[3]);
  assign or_108_nl = (mux_6_tmp[2:1]!=2'b11) | (mux_5_tmp[1:0]!=2'b00);
  assign mux_63_nl = MUX_s_1_2_2(or_108_nl, or_85_cse, mux_7_tmp[1]);
  assign mux_65_nl = MUX_s_1_2_2(mux_tmp_34, mux_63_nl, mux_7_tmp[0]);
  assign or_113_nl = (mux_6_tmp[3]) | mux_65_nl;
  assign mux_68_nl = MUX_s_1_2_2(mux_67_nl, or_113_nl, mux_6_tmp[0]);
  assign mux_69_nl = MUX_s_1_2_2(or_81_cse, mux_68_nl, mux_7_tmp[2]);
  assign and_dcpl_38 = (~ mux_69_nl) & and_dcpl_26 & and_dcpl_22;
  assign and_dcpl_39 = ~((mux_7_tmp[6:5]!=2'b00));
  assign and_dcpl_41 = ~((mux_7_tmp[4:3]!=2'b00));
  assign and_dcpl_42 = ~((mux_6_tmp[6:5]!=2'b00));
  assign and_dcpl_45 = ~((mux_5_tmp[6:5]!=2'b00));
  assign and_dcpl_47 = ~((mux_5_tmp[4:3]!=2'b00));
  assign and_dcpl_48 = (~ (mux_4_tmp[6])) & (mux_5_tmp[2]);
  assign not_tmp_66 = ~((mux_6_tmp[0]) & (mux_5_tmp[0]));
  assign or_125_nl = (mux_6_tmp[0]) | (~ (mux_5_tmp[0]));
  assign mux_74_nl = MUX_s_1_2_2(not_tmp_66, or_125_nl, mux_7_tmp[0]);
  assign nand_12_nl = ~((mux_7_tmp[1]) & (~ mux_74_nl));
  assign mux_71_nl = MUX_s_1_2_2((~ (mux_5_tmp[0])), (mux_5_tmp[0]), mux_6_tmp[0]);
  assign mux_72_nl = MUX_s_1_2_2(not_tmp_66, mux_71_nl, mux_7_tmp[0]);
  assign or_124_nl = (mux_7_tmp[0]) | (mux_6_tmp[0]) | (mux_5_tmp[0]);
  assign mux_73_nl = MUX_s_1_2_2(mux_72_nl, or_124_nl, mux_7_tmp[1]);
  assign mux_75_nl = MUX_s_1_2_2(nand_12_nl, mux_73_nl, mux_6_tmp[1]);
  assign and_148_nl = (mux_6_tmp[2]) & (mux_7_tmp[2]) & (~ mux_75_nl);
  assign or_122_nl = (mux_6_tmp[1]) | (mux_7_tmp[1:0]!=2'b11) | (mux_6_tmp[0]) |
      (~ (mux_5_tmp[0]));
  assign or_120_nl = (mux_6_tmp[1]) | (mux_7_tmp[1:0]!=2'b00) | (mux_6_tmp[0]) |
      (mux_5_tmp[0]);
  assign mux_70_nl = MUX_s_1_2_2(or_122_nl, or_120_nl, mux_7_tmp[2]);
  assign nor_34_nl = ~((mux_6_tmp[2]) | mux_70_nl);
  assign mux_76_nl = MUX_s_1_2_2(and_148_nl, nor_34_nl, mux_6_tmp[3]);
  assign and_dcpl_55 = mux_76_nl & and_dcpl_25 & and_dcpl_23 & (~ (mux_4_tmp[5]))
      & and_dcpl_48 & and_dcpl_47 & and_dcpl_45 & (~ (mux_6_tmp[4])) & and_dcpl_42
      & and_dcpl_41 & and_dcpl_39 & (~ (mux_5_tmp[1]));
  assign and_dcpl_58 = and_dcpl_12 & and_dcpl_10;
  assign and_dcpl_60 = ~((mux_5_tmp[6]) | (mux_6_tmp[4]));
  assign and_dcpl_63 = and_dcpl_18 & and_dcpl_16 & and_dcpl_60 & (~ (mux_6_tmp[5]));
  assign and_dcpl_64 = and_dcpl_63 & and_dcpl_58 & (~((mux_7_tmp[6]) | (mux_5_tmp[1])))
      & (mux_7_tmp[2]);
  assign and_dcpl_65 = ~((mux_4_tmp[5:4]!=2'b00));
  assign and_dcpl_69 = and_dcpl_24 & (mux_4_tmp[3:2]==2'b00) & and_dcpl_65 & (~ (mux_4_tmp[6]));
  assign or_tmp_75 = (mux_7_tmp[1]) | (mux_6_tmp[3:1]!=3'b011) | (mux_5_tmp[0]);
  assign nand_34_nl = ~((mux_6_tmp[3:1]==3'b011) & (mux_5_tmp[0]));
  assign or_130_nl = (mux_6_tmp[3:1]!=3'b010) | (~ (mux_5_tmp[0]));
  assign mux_tmp_63 = MUX_s_1_2_2(nand_34_nl, or_130_nl, mux_7_tmp[1]);
  assign or_134_nl = (mux_6_tmp[3:1]!=3'b100) | (mux_5_tmp[0]);
  assign or_133_nl = (mux_6_tmp[3:1]!=3'b011) | (mux_5_tmp[0]);
  assign mux_tmp_65 = MUX_s_1_2_2(or_134_nl, or_133_nl, mux_7_tmp[1]);
  assign mux_tmp_66 = MUX_s_1_2_2(mux_tmp_65, mux_tmp_63, mux_7_tmp[0]);
  assign mux_78_nl = MUX_s_1_2_2(mux_tmp_63, or_tmp_75, mux_7_tmp[0]);
  assign mux_81_nl = MUX_s_1_2_2(mux_tmp_66, mux_78_nl, mux_6_tmp[0]);
  assign and_dcpl_71 = (~ mux_81_nl) & and_dcpl_69 & and_dcpl_64;
  assign or_tmp_83 = (~ (mux_7_tmp[1])) | (mux_6_tmp[3:1]!=3'b010) | (~ (mux_5_tmp[0]));
  assign mux_tmp_68 = MUX_s_1_2_2(or_tmp_83, or_tmp_75, mux_7_tmp[0]);
  assign mux_83_nl = MUX_s_1_2_2(mux_tmp_66, mux_tmp_68, mux_6_tmp[0]);
  assign and_dcpl_73 = (~ mux_83_nl) & and_dcpl_69 & and_dcpl_64;
  assign mux_tmp_70 = MUX_s_1_2_2(mux_tmp_65, or_tmp_83, mux_7_tmp[0]);
  assign mux_85_nl = MUX_s_1_2_2(mux_tmp_70, mux_tmp_68, mux_6_tmp[0]);
  assign and_dcpl_75 = (~ mux_85_nl) & and_dcpl_69 & and_dcpl_64;
  assign or_143_nl = (mux_7_tmp[1:0]!=2'b01) | (mux_6_tmp[3:1]!=3'b011) | (mux_5_tmp[0]);
  assign mux_86_nl = MUX_s_1_2_2(mux_tmp_70, or_143_nl, mux_6_tmp[0]);
  assign and_dcpl_77 = (~ mux_86_nl) & and_dcpl_69 & and_dcpl_64;
  assign and_dcpl_87 = ~((mux_4_tmp[2:1]!=2'b00));
  assign or_149_nl = (mux_6_tmp[3:1]!=3'b100);
  assign or_147_nl = (mux_6_tmp[3:1]!=3'b011);
  assign mux_87_nl = MUX_s_1_2_2(or_149_nl, or_147_nl, mux_7_tmp[1]);
  assign or_1530_nl = (mux_7_tmp[0]) | mux_87_nl;
  assign or_1531_nl = (mux_7_tmp[1:0]!=2'b01) | (mux_6_tmp[3:1]!=3'b011);
  assign mux_88_nl = MUX_s_1_2_2(or_1530_nl, or_1531_nl, mux_6_tmp[0]);
  assign and_dcpl_92 = (~(mux_88_nl | (mux_4_tmp[0]))) & and_dcpl_87 & and_dcpl_23
      & and_dcpl_19 & (mux_5_tmp[2]) & and_dcpl_47 & and_dcpl_45 & and_dcpl_13 &
      (~ (mux_6_tmp[6])) & and_dcpl_41 & and_dcpl_39 & nor_25_cse & (mux_7_tmp[2]);
  assign and_dcpl_96 = ~((mux_7_tmp[6]) | (mux_5_tmp[0]));
  assign or_1532_nl = (mux_7_tmp[1:0]!=2'b10);
  assign or_1533_nl = (mux_7_tmp[1:0]!=2'b01);
  assign mux_89_nl = MUX_s_1_2_2(or_1532_nl, or_1533_nl, mux_6_tmp[0]);
  assign and_dcpl_110 = (~(mux_89_nl | (mux_4_tmp[0]))) & and_dcpl_87 & (~ (mux_4_tmp[3]))
      & and_dcpl_65 & and_dcpl_48 & and_dcpl_47 & (~ (mux_5_tmp[5])) & and_dcpl_60
      & and_dcpl_42 & and_dcpl_41 & (~ (mux_7_tmp[5])) & and_dcpl_96 & (~ (mux_5_tmp[1]))
      & (mux_7_tmp[2]) & (mux_6_tmp[3:1]==3'b011);
  assign and_dcpl_121 = and_dcpl_69 & and_dcpl_63 & and_dcpl_58 & and_dcpl_96 & (~
      (mux_5_tmp[1])) & (mux_7_tmp[2]) & (mux_6_tmp[3:1]==3'b011) & (mux_7_tmp[1:0]==2'b10)
      & (~ (mux_6_tmp[0]));
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      v_n_obs_sva <= 7'b0000000;
    end
    else if ( ((n_sva[2:0]==3'b111)) | and_149_cse ) begin
      v_n_obs_sva <= MUX_v_7_2_2(7'b0000000, v_n_obs_sva_dfm_1_mx0, unequal_tmp_3);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      run_sva <= 7'b0000000;
      reg_epsilon_triosy_obj_ld_cse <= 1'b0;
      is_random_rsci_idat <= 1'b0;
      valid_rsci_idat <= 1'b0;
      n_sva <= 7'b0000000;
    end
    else begin
      run_sva <= run_sva_2 & ({{6{epsilon_rsci_idat}}, epsilon_rsci_idat}) & ({{6{unequal_tmp_3}},
          unequal_tmp_3});
      reg_epsilon_triosy_obj_ld_cse <= 1'b1;
      is_random_rsci_idat <= ~((~((~((nu_3_sva_dfm_1_mx1!=7'b0000000) | (~ if_2_oif_472_land_1_lpi_1_dfm_mx0)))
          | if_2_lor_471_lpi_1_dfm_1_mx0)) | unequal_tmp_2);
      valid_rsci_idat <= ~ unequal_tmp_2;
      n_sva <= acc_tmp;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      nu_0_sva <= 7'b0000000;
    end
    else if ( (and_178_cse | mux_93_nl) & (n_sva[2:0]==3'b111) ) begin
      nu_0_sva <= MUX_v_7_2_2(7'b0000000, asn_25_mx0w1, unequal_tmp_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      nu_1_sva <= 7'b0000000;
    end
    else if ( (and_178_cse | mux_94_nl) & (n_sva[2:0]==3'b111) ) begin
      nu_1_sva <= MUX_v_7_2_2(7'b0000000, asn_24_mx0w0, unequal_tmp_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      nu_2_sva <= 7'b0000000;
    end
    else if ( (and_178_cse | mux_95_nl) & (n_sva[2:0]==3'b111) ) begin
      nu_2_sva <= MUX_v_7_2_2(7'b0000000, asn_22_mx0w0, unequal_tmp_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      nu_3_sva <= 7'b0000000;
    end
    else if ( (and_178_cse | mux_96_nl) & (n_sva[2:0]==3'b111) ) begin
      nu_3_sva <= MUX_v_7_2_2(7'b0000000, nu_3_sva_dfm_1_mx1, unequal_tmp_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_472_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( (n_sva[3:0]==4'b1111) & (~ if_2_if_if_2_if_or_471_tmp) & (n_sva[6:4]==3'b111)
        ) begin
      if_2_oif_472_land_1_lpi_1_dfm <= if_2_oif_472_land_1_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_lor_471_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ((acc_tmp!=7'b1111111)) & (n_sva==7'b1111111) ) begin
      if_2_lor_471_lpi_1_dfm_1 <= if_2_lor_471_lpi_1_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_14_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_28 | or_dcpl_38) ) begin
      if_2_oif_14_land_1_lpi_1_dfm <= if_2_oif_14_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_13_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_30 | or_dcpl_38) ) begin
      if_2_oif_13_land_1_lpi_1_dfm <= if_2_oif_13_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_12_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_32 | or_dcpl_38) ) begin
      if_2_oif_12_land_1_lpi_1_dfm <= if_2_oif_12_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_11_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_34 | or_dcpl_38) ) begin
      if_2_oif_11_land_1_lpi_1_dfm <= if_2_oif_11_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_10_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_36 | or_dcpl_38) ) begin
      if_2_oif_10_land_1_lpi_1_dfm <= if_2_oif_10_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_9_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_38 | or_dcpl_38) ) begin
      if_2_oif_9_land_1_lpi_1_dfm <= if_2_oif_9_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_8_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_55 | or_dcpl_38) ) begin
      if_2_oif_8_land_1_lpi_1_dfm <= if_2_oif_8_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_7_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_71 | or_dcpl_38) ) begin
      if_2_oif_7_land_1_lpi_1_dfm <= if_2_oif_7_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_6_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_73 | or_dcpl_38) ) begin
      if_2_oif_6_land_1_lpi_1_dfm <= if_2_oif_6_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_5_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_75 | or_dcpl_38) ) begin
      if_2_oif_5_land_1_lpi_1_dfm <= if_2_oif_5_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_4_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_77 | or_dcpl_38) ) begin
      if_2_oif_4_land_1_lpi_1_dfm <= if_2_oif_4_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_3_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_92 | or_dcpl_38) ) begin
      if_2_oif_3_land_1_lpi_1_dfm <= if_2_oif_3_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_2_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_110 | or_dcpl_38) ) begin
      if_2_oif_2_land_1_lpi_1_dfm <= if_2_oif_2_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_2_oif_1_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( ~(and_dcpl_121 | or_dcpl_38) ) begin
      if_2_oif_1_land_1_lpi_1_dfm <= if_2_oif_1_land_1_lpi_1_dfm_mx0w0;
    end
  end
  assign nor_56_nl = ~((v_n_obs_sva[6:1]!=6'b000000));
  assign nor_57_nl = ~((run_sva_2[6:1]!=6'b000000));
  assign mux_93_nl = MUX_s_1_2_2(nor_56_nl, nor_57_nl, and_149_cse);
  assign nor_58_nl = ~((v_n_obs_sva!=7'b0000010));
  assign nor_59_nl = ~((run_sva_2!=7'b0000010));
  assign mux_94_nl = MUX_s_1_2_2(nor_58_nl, nor_59_nl, and_149_cse);
  assign nor_60_nl = ~((v_n_obs_sva!=7'b0000011));
  assign nor_61_nl = ~((run_sva_2!=7'b0000011));
  assign mux_95_nl = MUX_s_1_2_2(nor_60_nl, nor_61_nl, and_149_cse);
  assign or_1545_nl = (v_n_obs_sva[6:2]!=5'b00000);
  assign or_1544_nl = (run_sva_2[6:2]!=5'b00000);
  assign mux_96_nl = MUX_s_1_2_2(or_1545_nl, or_1544_nl, and_149_cse);

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction

endmodule