magic
tech sky130A
magscale 1 2
timestamp 1713067979
<< nwell >>
rect -683 -384 683 384
<< pmos >>
rect -487 -164 -287 236
rect -229 -164 -29 236
rect 29 -164 229 236
rect 287 -164 487 236
<< pdiff >>
rect -545 224 -487 236
rect -545 -152 -533 224
rect -499 -152 -487 224
rect -545 -164 -487 -152
rect -287 224 -229 236
rect -287 -152 -275 224
rect -241 -152 -229 224
rect -287 -164 -229 -152
rect -29 224 29 236
rect -29 -152 -17 224
rect 17 -152 29 224
rect -29 -164 29 -152
rect 229 224 287 236
rect 229 -152 241 224
rect 275 -152 287 224
rect 229 -164 287 -152
rect 487 224 545 236
rect 487 -152 499 224
rect 533 -152 545 224
rect 487 -164 545 -152
<< pdiffc >>
rect -533 -152 -499 224
rect -275 -152 -241 224
rect -17 -152 17 224
rect 241 -152 275 224
rect 499 -152 533 224
<< nsubdiff >>
rect -647 314 -551 348
rect 551 314 647 348
rect -647 -314 -613 314
rect 613 -314 647 314
rect -647 -348 647 -314
<< nsubdiffcont >>
rect -551 314 551 348
<< poly >>
rect -487 236 -287 262
rect -229 236 -29 262
rect 29 236 229 262
rect 287 236 487 262
rect -487 -211 -287 -164
rect -487 -245 -471 -211
rect -303 -245 -287 -211
rect -487 -261 -287 -245
rect -229 -211 -29 -164
rect -229 -245 -213 -211
rect -45 -245 -29 -211
rect -229 -261 -29 -245
rect 29 -211 229 -164
rect 29 -245 45 -211
rect 213 -245 229 -211
rect 29 -261 229 -245
rect 287 -211 487 -164
rect 287 -245 303 -211
rect 471 -245 487 -211
rect 287 -261 487 -245
<< polycont >>
rect -471 -245 -303 -211
rect -213 -245 -45 -211
rect 45 -245 213 -211
rect 303 -245 471 -211
<< locali >>
rect -647 -314 -613 348
rect -533 224 -499 240
rect -533 -168 -499 -152
rect -275 224 -241 240
rect -275 -168 -241 -152
rect -17 224 17 240
rect -17 -168 17 -152
rect 241 224 275 240
rect 241 -168 275 -152
rect 499 224 533 240
rect 499 -168 533 -152
rect -487 -245 -471 -211
rect -303 -245 -287 -211
rect -229 -245 -213 -211
rect -45 -245 -29 -211
rect 29 -245 45 -211
rect 213 -245 229 -211
rect 287 -245 303 -211
rect 471 -245 487 -211
rect 613 -314 647 348
rect -647 -348 647 -314
<< viali >>
rect -613 314 -551 348
rect -551 314 551 348
rect 551 314 613 348
rect -533 -135 -499 15
rect -275 57 -241 207
rect -17 -135 17 15
rect 241 57 275 207
rect 499 -135 533 15
rect -471 -245 -303 -211
rect -213 -245 -45 -211
rect 45 -245 213 -211
rect 303 -245 471 -211
<< metal1 >>
rect -625 348 625 354
rect -625 314 -613 348
rect 613 314 625 348
rect -625 308 625 314
rect -281 207 -235 219
rect -281 57 -275 207
rect -241 57 -235 207
rect -281 45 -235 57
rect 235 207 281 219
rect 235 57 241 207
rect 275 57 281 207
rect 235 45 281 57
rect -539 15 -493 27
rect -539 -135 -533 15
rect -499 -135 -493 15
rect -539 -147 -493 -135
rect -23 15 23 27
rect -23 -135 -17 15
rect 17 -135 23 15
rect -23 -147 23 -135
rect 493 15 539 27
rect 493 -135 499 15
rect 533 -135 539 15
rect 493 -147 539 -135
rect -483 -211 -291 -205
rect -483 -245 -471 -211
rect -303 -245 -291 -211
rect -483 -251 -291 -245
rect -225 -211 -33 -205
rect -225 -245 -213 -211
rect -45 -245 -33 -211
rect -225 -251 -33 -245
rect 33 -211 225 -205
rect 33 -245 45 -211
rect 213 -245 225 -211
rect 33 -251 225 -245
rect 291 -211 483 -205
rect 291 -245 303 -211
rect 471 -245 483 -211
rect 291 -251 483 -245
<< properties >>
string FIXED_BBOX -630 -331 630 331
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
