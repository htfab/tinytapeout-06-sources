magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -1199 -379 1199 379
<< nmos >>
rect -1003 -169 -803 231
rect -745 -169 -545 231
rect -487 -169 -287 231
rect -229 -169 -29 231
rect 29 -169 229 231
rect 287 -169 487 231
rect 545 -169 745 231
rect 803 -169 1003 231
<< ndiff >>
rect -1061 219 -1003 231
rect -1061 -157 -1049 219
rect -1015 -157 -1003 219
rect -1061 -169 -1003 -157
rect -803 219 -745 231
rect -803 -157 -791 219
rect -757 -157 -745 219
rect -803 -169 -745 -157
rect -545 219 -487 231
rect -545 -157 -533 219
rect -499 -157 -487 219
rect -545 -169 -487 -157
rect -287 219 -229 231
rect -287 -157 -275 219
rect -241 -157 -229 219
rect -287 -169 -229 -157
rect -29 219 29 231
rect -29 -157 -17 219
rect 17 -157 29 219
rect -29 -169 29 -157
rect 229 219 287 231
rect 229 -157 241 219
rect 275 -157 287 219
rect 229 -169 287 -157
rect 487 219 545 231
rect 487 -157 499 219
rect 533 -157 545 219
rect 487 -169 545 -157
rect 745 219 803 231
rect 745 -157 757 219
rect 791 -157 803 219
rect 745 -169 803 -157
rect 1003 219 1061 231
rect 1003 -157 1015 219
rect 1049 -157 1061 219
rect 1003 -169 1061 -157
<< ndiffc >>
rect -1049 -157 -1015 219
rect -791 -157 -757 219
rect -533 -157 -499 219
rect -275 -157 -241 219
rect -17 -157 17 219
rect 241 -157 275 219
rect 499 -157 533 219
rect 757 -157 791 219
rect 1015 -157 1049 219
<< psubdiff >>
rect -1163 309 -1067 343
rect 1067 309 1163 343
rect -1163 247 -1129 309
rect 1129 247 1163 309
rect -1163 -309 -1129 -247
rect 1129 -309 1163 -247
rect -1163 -343 1163 -309
<< psubdiffcont >>
rect -1067 309 1067 343
rect -1163 -247 -1129 247
rect 1129 -247 1163 247
<< poly >>
rect -1003 231 -803 257
rect -745 231 -545 257
rect -487 231 -287 257
rect -229 231 -29 257
rect 29 231 229 257
rect 287 231 487 257
rect 545 231 745 257
rect 803 231 1003 257
rect -1003 -207 -803 -169
rect -1003 -241 -987 -207
rect -819 -241 -803 -207
rect -1003 -257 -803 -241
rect -745 -207 -545 -169
rect -745 -241 -729 -207
rect -561 -241 -545 -207
rect -745 -257 -545 -241
rect -487 -207 -287 -169
rect -487 -241 -471 -207
rect -303 -241 -287 -207
rect -487 -257 -287 -241
rect -229 -207 -29 -169
rect -229 -241 -213 -207
rect -45 -241 -29 -207
rect -229 -257 -29 -241
rect 29 -207 229 -169
rect 29 -241 45 -207
rect 213 -241 229 -207
rect 29 -257 229 -241
rect 287 -207 487 -169
rect 287 -241 303 -207
rect 471 -241 487 -207
rect 287 -257 487 -241
rect 545 -207 745 -169
rect 545 -241 561 -207
rect 729 -241 745 -207
rect 545 -257 745 -241
rect 803 -207 1003 -169
rect 803 -241 819 -207
rect 987 -241 1003 -207
rect 803 -257 1003 -241
<< polycont >>
rect -987 -241 -819 -207
rect -729 -241 -561 -207
rect -471 -241 -303 -207
rect -213 -241 -45 -207
rect 45 -241 213 -207
rect 303 -241 471 -207
rect 561 -241 729 -207
rect 819 -241 987 -207
<< locali >>
rect -1163 247 -1129 343
rect 1129 247 1163 343
rect -1049 219 -1015 235
rect -1049 -173 -1015 -157
rect -791 219 -757 235
rect -791 -173 -757 -157
rect -533 219 -499 235
rect -533 -173 -499 -157
rect -275 219 -241 235
rect -275 -173 -241 -157
rect -17 219 17 235
rect -17 -173 17 -157
rect 241 219 275 235
rect 241 -173 275 -157
rect 499 219 533 235
rect 499 -173 533 -157
rect 757 219 791 235
rect 757 -173 791 -157
rect 1015 219 1049 235
rect 1015 -173 1049 -157
rect -1003 -241 -987 -207
rect -819 -241 -803 -207
rect -745 -241 -729 -207
rect -561 -241 -545 -207
rect -487 -241 -471 -207
rect -303 -241 -287 -207
rect -229 -241 -213 -207
rect -45 -241 -29 -207
rect 29 -241 45 -207
rect 213 -241 229 -207
rect 287 -241 303 -207
rect 471 -241 487 -207
rect 545 -241 561 -207
rect 729 -241 745 -207
rect 803 -241 819 -207
rect 987 -241 1003 -207
rect -1163 -343 1163 -309
<< viali >>
rect -1129 309 -1067 343
rect -1067 309 1067 343
rect 1067 309 1129 343
rect -1163 -247 -1129 -62
rect -1049 52 -1015 202
rect -791 -140 -757 10
rect -533 52 -499 202
rect -275 -140 -241 10
rect -17 52 17 202
rect 241 -140 275 10
rect 499 52 533 202
rect 757 -140 791 10
rect 1015 52 1049 202
rect -987 -241 -819 -207
rect -729 -241 -561 -207
rect -471 -241 -303 -207
rect -213 -241 -45 -207
rect 45 -241 213 -207
rect 303 -241 471 -207
rect 561 -241 729 -207
rect 819 -241 987 -207
rect -1163 -309 -1129 -247
rect 1129 -247 1163 -62
rect 1129 -309 1163 -247
<< metal1 >>
rect -1141 343 1141 349
rect -1141 309 -1129 343
rect 1129 309 1141 343
rect -1141 303 1141 309
rect -1055 202 -1009 214
rect -1055 52 -1049 202
rect -1015 52 -1009 202
rect -1055 40 -1009 52
rect -539 202 -493 214
rect -539 52 -533 202
rect -499 52 -493 202
rect -539 40 -493 52
rect -23 202 23 214
rect -23 52 -17 202
rect 17 52 23 202
rect -23 40 23 52
rect 493 202 539 214
rect 493 52 499 202
rect 533 52 539 202
rect 493 40 539 52
rect 1009 202 1055 214
rect 1009 52 1015 202
rect 1049 52 1055 202
rect 1009 40 1055 52
rect -797 10 -751 22
rect -1169 -62 -1123 -50
rect -1169 -309 -1163 -62
rect -1129 -309 -1123 -62
rect -797 -140 -791 10
rect -757 -140 -751 10
rect -797 -152 -751 -140
rect -281 10 -235 22
rect -281 -140 -275 10
rect -241 -140 -235 10
rect -281 -152 -235 -140
rect 235 10 281 22
rect 235 -140 241 10
rect 275 -140 281 10
rect 235 -152 281 -140
rect 751 10 797 22
rect 751 -140 757 10
rect 791 -140 797 10
rect 751 -152 797 -140
rect 1123 -62 1169 -50
rect -999 -207 -807 -201
rect -999 -241 -987 -207
rect -819 -241 -807 -207
rect -999 -247 -807 -241
rect -741 -207 -549 -201
rect -741 -241 -729 -207
rect -561 -241 -549 -207
rect -741 -247 -549 -241
rect -483 -207 -291 -201
rect -483 -241 -471 -207
rect -303 -241 -291 -207
rect -483 -247 -291 -241
rect -225 -207 -33 -201
rect -225 -241 -213 -207
rect -45 -241 -33 -207
rect -225 -247 -33 -241
rect 33 -207 225 -201
rect 33 -241 45 -207
rect 213 -241 225 -207
rect 33 -247 225 -241
rect 291 -207 483 -201
rect 291 -241 303 -207
rect 471 -241 483 -207
rect 291 -247 483 -241
rect 549 -207 741 -201
rect 549 -241 561 -207
rect 729 -241 741 -207
rect 549 -247 741 -241
rect 807 -207 999 -201
rect 807 -241 819 -207
rect 987 -241 999 -207
rect 807 -247 999 -241
rect -1169 -321 -1123 -309
rect 1123 -309 1129 -62
rect 1163 -309 1169 -62
rect 1123 -321 1169 -309
<< properties >>
string FIXED_BBOX -1146 -326 1146 326
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
