magic
tech sky130A
magscale 1 2
timestamp 1713551876
<< metal1 >>
rect 19004 11954 21138 12054
rect 10962 11860 15460 11942
rect 10962 11004 11068 11860
rect 15322 11250 15460 11860
rect 15322 11004 15470 11250
rect 10962 10078 15470 11004
rect 19004 11018 19080 11954
rect 21044 11018 21138 11954
rect 19004 10132 21138 11018
rect 23416 11674 26996 11726
rect 23416 10966 23462 11674
rect 26906 10966 26996 11674
rect 23416 10178 26996 10966
rect 21397 8694 21743 8700
rect 20817 8348 21397 8694
rect 21397 8342 21743 8348
rect 10968 3648 16968 4786
rect 10968 2280 11078 3648
rect 12838 3624 16968 3648
rect 12838 2280 14866 3624
rect 10968 2256 14866 2280
rect 16736 2256 16968 3624
rect 10968 2134 16968 2256
rect 18860 3640 21256 7088
rect 25532 4618 29374 4622
rect 18860 2334 18928 3640
rect 21146 2334 21256 3640
rect 23420 3722 29374 4618
rect 23420 2624 23464 3722
rect 25520 3680 29374 3722
rect 25520 2704 27196 3680
rect 29232 2704 29374 3680
rect 25520 2624 29374 2704
rect 23420 2590 29374 2624
rect 23420 2588 25584 2590
rect 18860 2198 21256 2334
<< via1 >>
rect 11068 11004 15322 11860
rect 19080 11018 21044 11954
rect 23462 10966 26906 11674
rect 21397 8348 21743 8694
rect 11078 2280 12838 3648
rect 14866 2256 16736 3624
rect 18928 2334 21146 3640
rect 23464 2624 25520 3722
rect 27196 2704 29232 3680
<< metal2 >>
rect 25381 44776 25390 44778
rect 11549 44742 11558 44744
rect 2978 44686 11558 44742
rect 2978 43232 3034 44686
rect 11549 44684 11558 44686
rect 11618 44684 11627 44744
rect 19170 44720 25390 44776
rect 14776 44176 14836 44185
rect 9050 44118 14776 44174
rect 7024 43374 7084 43383
rect 7024 43305 7084 43314
rect 5000 43290 5060 43299
rect 5000 43221 5060 43230
rect 9050 43219 9106 44118
rect 14776 44107 14836 44116
rect 17135 43690 17144 43750
rect 17204 43690 17213 43750
rect 15907 43606 15916 43608
rect 15122 43550 15916 43606
rect 11063 43420 11072 43480
rect 11132 43420 11141 43480
rect 13823 43438 13832 43440
rect 11074 43366 11130 43420
rect 13098 43382 13832 43438
rect 13823 43380 13832 43382
rect 13892 43380 13901 43440
rect 15122 43380 15178 43550
rect 15907 43548 15916 43550
rect 15976 43548 15985 43608
rect 17146 43270 17202 43690
rect 9048 43210 9108 43219
rect 9048 43141 9108 43150
rect 9050 43138 9106 43141
rect 19170 43118 19226 44720
rect 25381 44718 25390 44720
rect 25450 44718 25459 44778
rect 28762 44284 28822 44293
rect 23218 44226 28762 44282
rect 21192 43628 21252 43637
rect 21192 43559 21252 43568
rect 21194 43350 21250 43559
rect 23218 43176 23274 44226
rect 28762 44215 28822 44224
rect 30238 44072 30298 44081
rect 30238 44003 30298 44012
rect 30240 43854 30296 44003
rect 27266 43798 30296 43854
rect 25240 43702 25300 43711
rect 25240 43633 25300 43642
rect 25242 43284 25298 43633
rect 27266 43304 27322 43798
rect 29279 43480 29288 43540
rect 29348 43480 29357 43540
rect 29290 43282 29346 43480
rect 19004 11954 21138 12054
rect 10986 11860 15414 11924
rect 10986 11004 11068 11860
rect 15322 11004 15414 11860
rect 10986 10940 15414 11004
rect 19004 11018 19080 11954
rect 21044 11018 21138 11954
rect 19004 10132 21138 11018
rect 23432 11674 26964 11700
rect 23432 10966 23462 11674
rect 26906 10966 26964 11674
rect 23432 10934 26964 10966
rect 21391 8348 21397 8694
rect 21743 8348 21749 8694
rect 16782 6190 18184 6310
rect 10398 5888 11182 6062
rect 10398 4363 10572 5888
rect 18064 4741 18184 6190
rect 21397 5968 21743 8348
rect 29228 6110 30226 6230
rect 21397 5966 22782 5968
rect 21397 5814 23612 5966
rect 21397 5810 22350 5814
rect 21445 5282 21619 5810
rect 21441 5118 21450 5282
rect 21614 5118 21623 5282
rect 21445 5113 21619 5118
rect 10398 4189 12003 4363
rect 12177 4189 12186 4363
rect 11030 3648 12972 3784
rect 11030 2280 11078 3648
rect 12838 2280 12972 3648
rect 11030 2170 12972 2280
rect 13346 1868 13466 4676
rect 13806 4544 14010 4664
rect 18060 4631 18069 4741
rect 18179 4631 18188 4741
rect 18064 4626 18184 4631
rect 12260 1748 13466 1868
rect 11287 1076 11397 1080
rect 12260 1076 12380 1748
rect 13890 1595 14010 4544
rect 14732 3624 16882 3770
rect 14732 2256 14866 3624
rect 16736 2256 16882 3624
rect 18870 3640 21196 3732
rect 18870 2334 18928 3640
rect 21146 2334 21196 3640
rect 23438 3722 25564 3772
rect 23438 2624 23464 3722
rect 25520 2624 25564 3722
rect 23438 2606 25564 2624
rect 18870 2290 21196 2334
rect 14732 2158 16882 2256
rect 13886 1485 13895 1595
rect 14005 1485 14014 1595
rect 13890 1480 14010 1485
rect 25794 1433 25914 4582
rect 26314 4122 26434 4572
rect 30106 4147 30226 6110
rect 26901 4122 27011 4126
rect 26314 4117 27016 4122
rect 26314 4007 26901 4117
rect 27011 4007 27016 4117
rect 30102 4037 30111 4147
rect 30221 4037 30230 4147
rect 30106 4032 30226 4037
rect 26314 4002 27016 4007
rect 26901 3998 27011 4002
rect 27168 3680 29272 3734
rect 27168 2704 27196 3680
rect 29232 2704 29272 3680
rect 27168 2678 29272 2704
rect 25790 1323 25799 1433
rect 25909 1323 25918 1433
rect 25794 1318 25914 1323
rect 11282 1071 12380 1076
rect 11282 961 11287 1071
rect 11397 961 12380 1071
rect 11282 956 12380 961
rect 11287 952 11397 956
<< via2 >>
rect 11558 44684 11618 44744
rect 7024 43314 7084 43374
rect 5000 43230 5060 43290
rect 14776 44116 14836 44176
rect 17144 43690 17204 43750
rect 11072 43420 11132 43480
rect 13832 43380 13892 43440
rect 15916 43548 15976 43608
rect 9048 43150 9108 43210
rect 25390 44718 25450 44778
rect 21192 43568 21252 43628
rect 28762 44224 28822 44284
rect 30238 44012 30298 44072
rect 25240 43642 25300 43702
rect 29288 43480 29348 43540
rect 11068 11004 15322 11860
rect 19080 11018 21044 11954
rect 23462 10966 26906 11674
rect 21450 5118 21614 5282
rect 12003 4189 12177 4363
rect 11078 2280 12838 3648
rect 18069 4631 18179 4741
rect 14866 2256 16736 3624
rect 18928 2334 21146 3640
rect 23464 2624 25520 3722
rect 13895 1485 14005 1595
rect 26901 4007 27011 4117
rect 30111 4037 30221 4147
rect 27196 2704 29232 3680
rect 25799 1323 25909 1433
rect 11287 961 11397 1071
<< metal3 >>
rect 11553 44744 11623 44749
rect 11998 44744 12004 44746
rect 11553 44684 11558 44744
rect 11618 44684 12004 44744
rect 11553 44679 11623 44684
rect 11998 44682 12004 44684
rect 12068 44682 12074 44746
rect 14990 44716 14996 44780
rect 15060 44716 15066 44780
rect 25385 44778 25455 44783
rect 25906 44778 25912 44780
rect 25385 44718 25390 44778
rect 25450 44718 25912 44778
rect 14044 44374 14108 44380
rect 7024 44312 14044 44372
rect 4998 43766 5062 43772
rect 4998 43696 5062 43702
rect 5000 43295 5060 43696
rect 7024 43379 7084 44312
rect 14044 44304 14108 44310
rect 14774 44366 14838 44372
rect 14774 44296 14838 44302
rect 14776 44181 14836 44296
rect 14771 44176 14841 44181
rect 14771 44116 14776 44176
rect 14836 44116 14841 44176
rect 14771 44111 14841 44116
rect 14998 43978 15058 44716
rect 25385 44713 25455 44718
rect 25906 44716 25912 44718
rect 25976 44716 25982 44780
rect 28760 44562 28824 44568
rect 28760 44492 28824 44498
rect 30236 44518 30300 44524
rect 28762 44289 28822 44492
rect 30236 44448 30300 44454
rect 28757 44284 28827 44289
rect 28757 44224 28762 44284
rect 28822 44224 28827 44284
rect 28757 44219 28827 44224
rect 30238 44077 30298 44448
rect 30233 44072 30303 44077
rect 12120 43918 15058 43978
rect 21190 44032 21254 44038
rect 30233 44012 30238 44072
rect 30298 44012 30303 44072
rect 30233 44007 30303 44012
rect 21190 43962 21254 43968
rect 11067 43480 11137 43485
rect 12120 43480 12180 43918
rect 17139 43750 17209 43755
rect 17430 43750 17436 43752
rect 17139 43690 17144 43750
rect 17204 43690 17436 43750
rect 17139 43685 17209 43690
rect 17430 43688 17436 43690
rect 17500 43688 17506 43752
rect 21192 43633 21252 43962
rect 25238 43916 25302 43922
rect 25238 43846 25302 43852
rect 25240 43707 25300 43846
rect 25235 43702 25305 43707
rect 25235 43642 25240 43702
rect 25300 43642 25305 43702
rect 25235 43637 25305 43642
rect 21187 43628 21257 43633
rect 15911 43608 15981 43613
rect 16762 43610 16826 43616
rect 15911 43548 15916 43608
rect 15976 43548 16762 43608
rect 15911 43543 15981 43548
rect 21187 43568 21192 43628
rect 21252 43568 21257 43628
rect 21187 43563 21257 43568
rect 16762 43540 16826 43546
rect 29283 43540 29353 43545
rect 30724 43540 30730 43542
rect 7019 43374 7089 43379
rect 7019 43314 7024 43374
rect 7084 43314 7089 43374
rect 7019 43309 7089 43314
rect 4995 43290 5065 43295
rect 4995 43230 5000 43290
rect 5060 43230 5065 43290
rect 4995 43225 5065 43230
rect 9048 43215 9108 43440
rect 11067 43420 11072 43480
rect 11132 43420 12180 43480
rect 29283 43480 29288 43540
rect 29348 43480 30730 43540
rect 29283 43475 29353 43480
rect 30724 43478 30730 43480
rect 30794 43478 30800 43542
rect 13827 43440 13897 43445
rect 14404 43442 14468 43448
rect 11067 43415 11137 43420
rect 13827 43380 13832 43440
rect 13892 43380 14404 43440
rect 13827 43375 13897 43380
rect 14404 43372 14468 43378
rect 9043 43210 9113 43215
rect 9043 43150 9048 43210
rect 9108 43150 9113 43210
rect 9043 43145 9113 43150
rect 5540 14854 5852 14856
rect 5526 14536 5536 14854
rect 5860 14536 5870 14854
rect 12506 14536 12516 14880
rect 12832 14536 12842 14880
rect 19478 14860 19790 14868
rect 5540 12626 5852 14536
rect 5540 12608 10766 12626
rect 12528 12616 12840 14536
rect 19468 14516 19478 14860
rect 19790 14516 19800 14860
rect 26464 14806 26776 14812
rect 5540 12196 10222 12608
rect 10736 12196 10766 12608
rect 12510 12226 12520 12616
rect 12836 12226 12846 12616
rect 19478 12608 19790 14516
rect 26464 14512 26482 14806
rect 26776 14512 26786 14806
rect 12528 12222 12840 12226
rect 19464 12218 19474 12608
rect 19790 12218 19800 12608
rect 26464 12554 26776 14512
rect 19478 12210 19790 12218
rect 5540 12174 10766 12196
rect 26434 12154 26444 12554
rect 26868 12154 26878 12554
rect 19004 11954 21138 12054
rect 10986 11860 15414 11924
rect 10986 11004 11068 11860
rect 15322 11004 15414 11860
rect 10986 10940 15414 11004
rect 19004 11018 19080 11954
rect 21044 11018 21138 11954
rect 19004 10132 21138 11018
rect 23432 11674 26964 11700
rect 23432 10966 23462 11674
rect 26906 10966 26964 11674
rect 23432 10934 26964 10966
rect 17449 5282 21619 5287
rect 17449 5118 21450 5282
rect 21614 5118 21619 5282
rect 17449 5113 21619 5118
rect 11998 4363 12182 4368
rect 17449 4363 17623 5113
rect 11998 4189 12003 4363
rect 12177 4189 17623 4363
rect 18064 4741 18184 4746
rect 18064 4631 18069 4741
rect 18179 4631 18184 4741
rect 11998 4184 12182 4189
rect 11030 3648 12972 3784
rect 11030 2280 11078 3648
rect 12838 2280 12972 3648
rect 11030 2170 12972 2280
rect 14732 3624 16882 3770
rect 14732 2256 14866 3624
rect 16736 2256 16882 3624
rect 14732 2158 16882 2256
rect 13648 1595 14010 1600
rect 13648 1485 13895 1595
rect 14005 1485 14010 1595
rect 13648 1480 14010 1485
rect 9233 1076 9351 1081
rect 9232 1075 11402 1076
rect 9232 957 9233 1075
rect 9351 1071 11402 1075
rect 9351 961 11287 1071
rect 11397 961 11402 1071
rect 9351 957 11402 961
rect 9232 956 11402 957
rect 9233 951 9351 956
rect 13648 567 13768 1480
rect 18064 585 18184 4631
rect 30106 4147 30226 4152
rect 26896 4117 27016 4122
rect 26896 4007 26901 4117
rect 27011 4007 27016 4117
rect 18870 3640 21196 3732
rect 18870 2334 18928 3640
rect 21146 2334 21196 3640
rect 23438 3722 25564 3772
rect 23438 2624 23464 3722
rect 25520 2624 25564 3722
rect 23438 2606 25564 2624
rect 18870 2290 21196 2334
rect 22480 1433 25914 1438
rect 22480 1323 25799 1433
rect 25909 1323 25914 1433
rect 22480 1318 25914 1323
rect 22480 627 22600 1318
rect 26896 673 27016 4007
rect 30106 4037 30111 4147
rect 30221 4037 30226 4147
rect 27168 3680 29272 3734
rect 27168 2704 27196 3680
rect 29232 2704 29272 3680
rect 27168 2678 29272 2704
rect 30106 941 30226 4037
rect 30101 823 30107 941
rect 30225 823 30231 941
rect 30106 822 30226 823
rect 13643 449 13649 567
rect 13767 449 13773 567
rect 18059 467 18065 585
rect 18183 467 18189 585
rect 22475 509 22481 627
rect 22599 509 22605 627
rect 26891 555 26897 673
rect 27015 555 27021 673
rect 30106 614 30226 620
rect 26896 554 27016 555
rect 22480 508 22600 509
rect 30101 495 30106 613
rect 30226 495 30231 613
rect 30106 488 30226 494
rect 18064 466 18184 467
rect 13648 448 13768 449
<< via3 >>
rect 12004 44682 12068 44746
rect 14996 44716 15060 44780
rect 4998 43702 5062 43766
rect 14044 44310 14108 44374
rect 14774 44302 14838 44366
rect 25912 44716 25976 44780
rect 28760 44498 28824 44562
rect 30236 44454 30300 44518
rect 21190 43968 21254 44032
rect 17436 43688 17500 43752
rect 25238 43852 25302 43916
rect 16762 43546 16826 43610
rect 30730 43478 30794 43542
rect 14404 43378 14468 43442
rect 5536 14536 5860 14854
rect 12516 14536 12832 14880
rect 19478 14516 19790 14860
rect 10222 12196 10736 12608
rect 12520 12226 12836 12616
rect 26482 14512 26776 14806
rect 19474 12218 19790 12608
rect 26444 12154 26868 12554
rect 11068 11004 15322 11860
rect 19080 11018 21044 11954
rect 23462 10966 26906 11674
rect 11078 2280 12838 3648
rect 14866 2256 16736 3624
rect 9233 957 9351 1075
rect 18928 2334 21146 3640
rect 23464 2624 25520 3722
rect 27196 2704 29232 3680
rect 30107 823 30225 941
rect 13649 449 13767 567
rect 18065 467 18183 585
rect 22481 509 22599 627
rect 26897 555 27015 673
rect 30106 494 30226 614
<< metal4 >>
rect 798 44878 858 45152
rect 1534 44878 1594 45152
rect 2270 44878 2330 45152
rect 3006 44878 3066 45152
rect 3742 44878 3802 45152
rect 4478 44878 4538 45152
rect 5214 44878 5274 45152
rect 5950 44878 6010 45152
rect 6686 44878 6746 45152
rect 7422 44878 7482 45152
rect 8158 44878 8218 45152
rect 8894 44878 8954 45152
rect 9630 44878 9690 45152
rect 10366 44878 10426 45152
rect 11102 44878 11162 45152
rect 11838 44878 11898 45152
rect 410 44818 11898 44878
rect 12574 45050 12634 45152
rect 12574 44831 12636 45050
rect 13310 44952 13370 45152
rect 410 44152 470 44818
rect 12573 44750 12636 44831
rect 13308 44842 13370 44952
rect 14046 44850 14106 45152
rect 13308 44754 13372 44842
rect 12003 44746 12069 44747
rect 12003 44682 12004 44746
rect 12068 44744 12069 44746
rect 12573 44745 12635 44750
rect 12267 44744 12635 44745
rect 12068 44684 12635 44744
rect 12068 44682 12069 44684
rect 12267 44683 12635 44684
rect 12003 44681 12069 44682
rect 13312 44534 13372 44754
rect 5000 44474 13372 44534
rect 14046 44754 14108 44850
rect 14782 44760 14842 45152
rect 200 14156 500 44152
rect 5000 43767 5060 44474
rect 14046 44375 14106 44754
rect 14776 44702 14842 44760
rect 14995 44780 15061 44781
rect 14995 44716 14996 44780
rect 15060 44778 15061 44780
rect 15518 44778 15578 45152
rect 15060 44718 15580 44778
rect 15060 44716 15061 44718
rect 14995 44715 15061 44716
rect 14043 44374 14109 44375
rect 14043 44310 14044 44374
rect 14108 44310 14109 44374
rect 14776 44367 14836 44702
rect 14043 44309 14109 44310
rect 14773 44366 14839 44367
rect 14773 44302 14774 44366
rect 14838 44302 14839 44366
rect 14773 44301 14839 44302
rect 16254 44102 16314 45152
rect 16990 44806 17050 45152
rect 17726 44898 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 16990 44674 17052 44806
rect 16992 44316 17052 44674
rect 16252 44004 16314 44102
rect 16764 44256 17052 44316
rect 17724 44674 17786 44898
rect 25911 44780 25977 44781
rect 25911 44716 25912 44780
rect 25976 44778 25977 44780
rect 27294 44778 27354 45152
rect 28030 45096 28090 45152
rect 25976 44718 27354 44778
rect 28026 44952 28090 45096
rect 28766 45070 28826 45152
rect 28762 44952 28826 45070
rect 29502 45028 29562 45152
rect 29496 44952 29562 45028
rect 25976 44716 25977 44718
rect 25911 44715 25977 44716
rect 16252 43866 16312 44004
rect 14560 43806 16312 43866
rect 4997 43766 5063 43767
rect 4997 43702 4998 43766
rect 5062 43702 5063 43766
rect 4997 43701 5063 43702
rect 14403 43442 14469 43443
rect 14403 43378 14404 43442
rect 14468 43440 14469 43442
rect 14560 43440 14620 43806
rect 16764 43611 16824 44256
rect 17435 43752 17501 43753
rect 17435 43688 17436 43752
rect 17500 43750 17501 43752
rect 17724 43750 17784 44674
rect 28026 44594 28086 44952
rect 21192 44534 28086 44594
rect 28762 44563 28822 44952
rect 28759 44562 28825 44563
rect 21192 44033 21252 44534
rect 28759 44498 28760 44562
rect 28824 44498 28825 44562
rect 28759 44497 28825 44498
rect 29496 44092 29556 44952
rect 30238 44519 30298 45152
rect 30235 44518 30301 44519
rect 30235 44454 30236 44518
rect 30300 44454 30301 44518
rect 30235 44453 30301 44454
rect 21189 44032 21255 44033
rect 21189 43968 21190 44032
rect 21254 43968 21255 44032
rect 21189 43967 21255 43968
rect 25240 44032 29556 44092
rect 25240 43917 25300 44032
rect 25237 43916 25303 43917
rect 25237 43852 25238 43916
rect 25302 43852 25303 43916
rect 25237 43851 25303 43852
rect 17500 43690 17784 43750
rect 17500 43688 17501 43690
rect 17435 43687 17501 43688
rect 16761 43610 16827 43611
rect 16761 43546 16762 43610
rect 16826 43546 16827 43610
rect 16761 43545 16827 43546
rect 30729 43542 30795 43543
rect 30729 43478 30730 43542
rect 30794 43540 30795 43542
rect 30974 43540 31034 45152
rect 31710 44952 31770 45152
rect 30794 43480 31034 43540
rect 30794 43478 30795 43480
rect 30729 43477 30795 43478
rect 14468 43380 14620 43440
rect 14468 43378 14469 43380
rect 14403 43377 14469 43378
rect 5536 14855 5876 15342
rect 5535 14854 5876 14855
rect 5535 14536 5536 14854
rect 5860 14536 5876 14854
rect 5535 14535 5861 14536
rect 9040 14156 9340 15264
rect 12516 14881 12838 15368
rect 12515 14880 12838 14881
rect 12515 14536 12516 14880
rect 12832 14536 12838 14880
rect 12515 14535 12833 14536
rect 16010 14156 16310 15350
rect 19478 14861 19816 15368
rect 19477 14860 19816 14861
rect 19477 14516 19478 14860
rect 19790 14516 19816 14860
rect 19477 14515 19791 14516
rect 22990 14156 23290 15156
rect 26450 14806 26788 15368
rect 26450 14512 26482 14806
rect 26776 14516 26788 14806
rect 26776 14512 26777 14516
rect 26481 14511 26777 14512
rect 29952 14156 30252 15592
rect 200 13856 30252 14156
rect 200 3796 500 13856
rect 29982 12624 31442 12630
rect 31616 12624 31916 44152
rect 10198 12616 31916 12624
rect 10198 12608 12520 12616
rect 10198 12196 10222 12608
rect 10736 12226 12520 12608
rect 12836 12608 31916 12616
rect 12836 12226 19474 12608
rect 10736 12218 19474 12226
rect 19790 12554 31916 12608
rect 19790 12218 26444 12554
rect 10736 12196 26444 12218
rect 10198 12154 26444 12196
rect 26868 12154 31916 12554
rect 10198 11954 31916 12154
rect 10198 11860 19080 11954
rect 10198 11004 11068 11860
rect 15322 11018 19080 11860
rect 21044 11674 31916 11954
rect 21044 11018 23462 11674
rect 15322 11004 23462 11018
rect 10198 10966 23462 11004
rect 26906 10966 31916 11674
rect 10198 10942 31916 10966
rect 10198 10918 18764 10942
rect 21574 10918 31916 10942
rect 29982 10914 31442 10918
rect 19922 3800 20160 3808
rect 10264 3796 30594 3800
rect 200 3722 30594 3796
rect 200 3648 23464 3722
rect 200 2280 11078 3648
rect 12838 3640 23464 3648
rect 12838 3624 18928 3640
rect 12838 2280 14866 3624
rect 200 2256 14866 2280
rect 16736 2334 18928 3624
rect 21146 2624 23464 3640
rect 25520 3680 30594 3722
rect 25520 2704 27196 3680
rect 29232 2704 30594 3680
rect 25520 2624 30594 2704
rect 21146 2334 30594 2624
rect 16736 2256 30594 2334
rect 200 2094 30594 2256
rect 200 1000 500 2094
rect 9232 1075 9352 1076
rect 9232 957 9233 1075
rect 9351 957 9352 1075
rect 31616 1000 31916 10918
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 957
rect 30106 941 30226 942
rect 30106 823 30107 941
rect 30225 823 30226 941
rect 26896 673 27016 674
rect 22480 627 22600 628
rect 18064 585 18184 586
rect 13648 567 13768 568
rect 13648 449 13649 567
rect 13767 449 13768 567
rect 13648 0 13768 449
rect 18064 467 18065 585
rect 18183 467 18184 585
rect 18064 0 18184 467
rect 22480 509 22481 627
rect 22599 509 22600 627
rect 22480 0 22600 509
rect 26896 555 26897 673
rect 27015 555 27016 673
rect 30106 615 30226 823
rect 26896 0 27016 555
rect 30105 614 30227 615
rect 30105 494 30106 614
rect 30226 494 31432 614
rect 30105 493 30227 494
rect 31312 0 31432 494
use opamp  opamp_0
timestamp 1713422843
transform 1 0 21426 0 1 7506
box 1988 -3100 7988 2900
use opamp  opamp_1
timestamp 1713422843
transform 1 0 8980 0 1 7586
box 1988 -3100 7988 2900
use top  top_0
timestamp 1713551075
transform 1 0 1672 0 1 14438
box 514 496 28587 29000
use vbias_resistor  vbias_resistor_0
timestamp 1713420874
transform 1 0 17820 0 1 7778
box 1048 -958 3482 2578
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 31616 1000 31916 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
