magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -2102 -719 2102 719
<< nmos >>
rect -1906 109 -1706 509
rect -1648 109 -1448 509
rect -1390 109 -1190 509
rect -1132 109 -932 509
rect -874 109 -674 509
rect -616 109 -416 509
rect -358 109 -158 509
rect -100 109 100 509
rect 158 109 358 509
rect 416 109 616 509
rect 674 109 874 509
rect 932 109 1132 509
rect 1190 109 1390 509
rect 1448 109 1648 509
rect 1706 109 1906 509
rect -1906 -509 -1706 -109
rect -1648 -509 -1448 -109
rect -1390 -509 -1190 -109
rect -1132 -509 -932 -109
rect -874 -509 -674 -109
rect -616 -509 -416 -109
rect -358 -509 -158 -109
rect -100 -509 100 -109
rect 158 -509 358 -109
rect 416 -509 616 -109
rect 674 -509 874 -109
rect 932 -509 1132 -109
rect 1190 -509 1390 -109
rect 1448 -509 1648 -109
rect 1706 -509 1906 -109
<< ndiff >>
rect -1964 497 -1906 509
rect -1964 121 -1952 497
rect -1918 121 -1906 497
rect -1964 109 -1906 121
rect -1706 497 -1648 509
rect -1706 121 -1694 497
rect -1660 121 -1648 497
rect -1706 109 -1648 121
rect -1448 497 -1390 509
rect -1448 121 -1436 497
rect -1402 121 -1390 497
rect -1448 109 -1390 121
rect -1190 497 -1132 509
rect -1190 121 -1178 497
rect -1144 121 -1132 497
rect -1190 109 -1132 121
rect -932 497 -874 509
rect -932 121 -920 497
rect -886 121 -874 497
rect -932 109 -874 121
rect -674 497 -616 509
rect -674 121 -662 497
rect -628 121 -616 497
rect -674 109 -616 121
rect -416 497 -358 509
rect -416 121 -404 497
rect -370 121 -358 497
rect -416 109 -358 121
rect -158 497 -100 509
rect -158 121 -146 497
rect -112 121 -100 497
rect -158 109 -100 121
rect 100 497 158 509
rect 100 121 112 497
rect 146 121 158 497
rect 100 109 158 121
rect 358 497 416 509
rect 358 121 370 497
rect 404 121 416 497
rect 358 109 416 121
rect 616 497 674 509
rect 616 121 628 497
rect 662 121 674 497
rect 616 109 674 121
rect 874 497 932 509
rect 874 121 886 497
rect 920 121 932 497
rect 874 109 932 121
rect 1132 497 1190 509
rect 1132 121 1144 497
rect 1178 121 1190 497
rect 1132 109 1190 121
rect 1390 497 1448 509
rect 1390 121 1402 497
rect 1436 121 1448 497
rect 1390 109 1448 121
rect 1648 497 1706 509
rect 1648 121 1660 497
rect 1694 121 1706 497
rect 1648 109 1706 121
rect 1906 497 1964 509
rect 1906 121 1918 497
rect 1952 121 1964 497
rect 1906 109 1964 121
rect -1964 -121 -1906 -109
rect -1964 -497 -1952 -121
rect -1918 -497 -1906 -121
rect -1964 -509 -1906 -497
rect -1706 -121 -1648 -109
rect -1706 -497 -1694 -121
rect -1660 -497 -1648 -121
rect -1706 -509 -1648 -497
rect -1448 -121 -1390 -109
rect -1448 -497 -1436 -121
rect -1402 -497 -1390 -121
rect -1448 -509 -1390 -497
rect -1190 -121 -1132 -109
rect -1190 -497 -1178 -121
rect -1144 -497 -1132 -121
rect -1190 -509 -1132 -497
rect -932 -121 -874 -109
rect -932 -497 -920 -121
rect -886 -497 -874 -121
rect -932 -509 -874 -497
rect -674 -121 -616 -109
rect -674 -497 -662 -121
rect -628 -497 -616 -121
rect -674 -509 -616 -497
rect -416 -121 -358 -109
rect -416 -497 -404 -121
rect -370 -497 -358 -121
rect -416 -509 -358 -497
rect -158 -121 -100 -109
rect -158 -497 -146 -121
rect -112 -497 -100 -121
rect -158 -509 -100 -497
rect 100 -121 158 -109
rect 100 -497 112 -121
rect 146 -497 158 -121
rect 100 -509 158 -497
rect 358 -121 416 -109
rect 358 -497 370 -121
rect 404 -497 416 -121
rect 358 -509 416 -497
rect 616 -121 674 -109
rect 616 -497 628 -121
rect 662 -497 674 -121
rect 616 -509 674 -497
rect 874 -121 932 -109
rect 874 -497 886 -121
rect 920 -497 932 -121
rect 874 -509 932 -497
rect 1132 -121 1190 -109
rect 1132 -497 1144 -121
rect 1178 -497 1190 -121
rect 1132 -509 1190 -497
rect 1390 -121 1448 -109
rect 1390 -497 1402 -121
rect 1436 -497 1448 -121
rect 1390 -509 1448 -497
rect 1648 -121 1706 -109
rect 1648 -497 1660 -121
rect 1694 -497 1706 -121
rect 1648 -509 1706 -497
rect 1906 -121 1964 -109
rect 1906 -497 1918 -121
rect 1952 -497 1964 -121
rect 1906 -509 1964 -497
<< ndiffc >>
rect -1952 121 -1918 497
rect -1694 121 -1660 497
rect -1436 121 -1402 497
rect -1178 121 -1144 497
rect -920 121 -886 497
rect -662 121 -628 497
rect -404 121 -370 497
rect -146 121 -112 497
rect 112 121 146 497
rect 370 121 404 497
rect 628 121 662 497
rect 886 121 920 497
rect 1144 121 1178 497
rect 1402 121 1436 497
rect 1660 121 1694 497
rect 1918 121 1952 497
rect -1952 -497 -1918 -121
rect -1694 -497 -1660 -121
rect -1436 -497 -1402 -121
rect -1178 -497 -1144 -121
rect -920 -497 -886 -121
rect -662 -497 -628 -121
rect -404 -497 -370 -121
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect 370 -497 404 -121
rect 628 -497 662 -121
rect 886 -497 920 -121
rect 1144 -497 1178 -121
rect 1402 -497 1436 -121
rect 1660 -497 1694 -121
rect 1918 -497 1952 -121
<< psubdiff >>
rect -2066 649 2066 683
rect -2066 587 -2032 649
rect 2032 587 2066 649
rect -2066 -649 -2032 -587
rect 2032 -649 2066 -587
rect -2066 -683 -1970 -649
rect 1970 -683 2066 -649
<< psubdiffcont >>
rect -2066 -587 -2032 587
rect 2032 -587 2066 587
rect -1970 -683 1970 -649
<< poly >>
rect -1906 581 -1706 597
rect -1906 547 -1890 581
rect -1722 547 -1706 581
rect -1906 509 -1706 547
rect -1648 581 -1448 597
rect -1648 547 -1632 581
rect -1464 547 -1448 581
rect -1648 509 -1448 547
rect -1390 581 -1190 597
rect -1390 547 -1374 581
rect -1206 547 -1190 581
rect -1390 509 -1190 547
rect -1132 581 -932 597
rect -1132 547 -1116 581
rect -948 547 -932 581
rect -1132 509 -932 547
rect -874 581 -674 597
rect -874 547 -858 581
rect -690 547 -674 581
rect -874 509 -674 547
rect -616 581 -416 597
rect -616 547 -600 581
rect -432 547 -416 581
rect -616 509 -416 547
rect -358 581 -158 597
rect -358 547 -342 581
rect -174 547 -158 581
rect -358 509 -158 547
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 509 100 547
rect 158 581 358 597
rect 158 547 174 581
rect 342 547 358 581
rect 158 509 358 547
rect 416 581 616 597
rect 416 547 432 581
rect 600 547 616 581
rect 416 509 616 547
rect 674 581 874 597
rect 674 547 690 581
rect 858 547 874 581
rect 674 509 874 547
rect 932 581 1132 597
rect 932 547 948 581
rect 1116 547 1132 581
rect 932 509 1132 547
rect 1190 581 1390 597
rect 1190 547 1206 581
rect 1374 547 1390 581
rect 1190 509 1390 547
rect 1448 581 1648 597
rect 1448 547 1464 581
rect 1632 547 1648 581
rect 1448 509 1648 547
rect 1706 581 1906 597
rect 1706 547 1722 581
rect 1890 547 1906 581
rect 1706 509 1906 547
rect -1906 71 -1706 109
rect -1906 37 -1890 71
rect -1722 37 -1706 71
rect -1906 21 -1706 37
rect -1648 71 -1448 109
rect -1648 37 -1632 71
rect -1464 37 -1448 71
rect -1648 21 -1448 37
rect -1390 71 -1190 109
rect -1390 37 -1374 71
rect -1206 37 -1190 71
rect -1390 21 -1190 37
rect -1132 71 -932 109
rect -1132 37 -1116 71
rect -948 37 -932 71
rect -1132 21 -932 37
rect -874 71 -674 109
rect -874 37 -858 71
rect -690 37 -674 71
rect -874 21 -674 37
rect -616 71 -416 109
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 109
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 109
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 109
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect 674 71 874 109
rect 674 37 690 71
rect 858 37 874 71
rect 674 21 874 37
rect 932 71 1132 109
rect 932 37 948 71
rect 1116 37 1132 71
rect 932 21 1132 37
rect 1190 71 1390 109
rect 1190 37 1206 71
rect 1374 37 1390 71
rect 1190 21 1390 37
rect 1448 71 1648 109
rect 1448 37 1464 71
rect 1632 37 1648 71
rect 1448 21 1648 37
rect 1706 71 1906 109
rect 1706 37 1722 71
rect 1890 37 1906 71
rect 1706 21 1906 37
rect -1906 -37 -1706 -21
rect -1906 -71 -1890 -37
rect -1722 -71 -1706 -37
rect -1906 -109 -1706 -71
rect -1648 -37 -1448 -21
rect -1648 -71 -1632 -37
rect -1464 -71 -1448 -37
rect -1648 -109 -1448 -71
rect -1390 -37 -1190 -21
rect -1390 -71 -1374 -37
rect -1206 -71 -1190 -37
rect -1390 -109 -1190 -71
rect -1132 -37 -932 -21
rect -1132 -71 -1116 -37
rect -948 -71 -932 -37
rect -1132 -109 -932 -71
rect -874 -37 -674 -21
rect -874 -71 -858 -37
rect -690 -71 -674 -37
rect -874 -109 -674 -71
rect -616 -37 -416 -21
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -616 -109 -416 -71
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -109 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -109 358 -71
rect 416 -37 616 -21
rect 416 -71 432 -37
rect 600 -71 616 -37
rect 416 -109 616 -71
rect 674 -37 874 -21
rect 674 -71 690 -37
rect 858 -71 874 -37
rect 674 -109 874 -71
rect 932 -37 1132 -21
rect 932 -71 948 -37
rect 1116 -71 1132 -37
rect 932 -109 1132 -71
rect 1190 -37 1390 -21
rect 1190 -71 1206 -37
rect 1374 -71 1390 -37
rect 1190 -109 1390 -71
rect 1448 -37 1648 -21
rect 1448 -71 1464 -37
rect 1632 -71 1648 -37
rect 1448 -109 1648 -71
rect 1706 -37 1906 -21
rect 1706 -71 1722 -37
rect 1890 -71 1906 -37
rect 1706 -109 1906 -71
rect -1906 -547 -1706 -509
rect -1906 -581 -1890 -547
rect -1722 -581 -1706 -547
rect -1906 -597 -1706 -581
rect -1648 -547 -1448 -509
rect -1648 -581 -1632 -547
rect -1464 -581 -1448 -547
rect -1648 -597 -1448 -581
rect -1390 -547 -1190 -509
rect -1390 -581 -1374 -547
rect -1206 -581 -1190 -547
rect -1390 -597 -1190 -581
rect -1132 -547 -932 -509
rect -1132 -581 -1116 -547
rect -948 -581 -932 -547
rect -1132 -597 -932 -581
rect -874 -547 -674 -509
rect -874 -581 -858 -547
rect -690 -581 -674 -547
rect -874 -597 -674 -581
rect -616 -547 -416 -509
rect -616 -581 -600 -547
rect -432 -581 -416 -547
rect -616 -597 -416 -581
rect -358 -547 -158 -509
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -358 -597 -158 -581
rect -100 -547 100 -509
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
rect 158 -547 358 -509
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 158 -597 358 -581
rect 416 -547 616 -509
rect 416 -581 432 -547
rect 600 -581 616 -547
rect 416 -597 616 -581
rect 674 -547 874 -509
rect 674 -581 690 -547
rect 858 -581 874 -547
rect 674 -597 874 -581
rect 932 -547 1132 -509
rect 932 -581 948 -547
rect 1116 -581 1132 -547
rect 932 -597 1132 -581
rect 1190 -547 1390 -509
rect 1190 -581 1206 -547
rect 1374 -581 1390 -547
rect 1190 -597 1390 -581
rect 1448 -547 1648 -509
rect 1448 -581 1464 -547
rect 1632 -581 1648 -547
rect 1448 -597 1648 -581
rect 1706 -547 1906 -509
rect 1706 -581 1722 -547
rect 1890 -581 1906 -547
rect 1706 -597 1906 -581
<< polycont >>
rect -1890 547 -1722 581
rect -1632 547 -1464 581
rect -1374 547 -1206 581
rect -1116 547 -948 581
rect -858 547 -690 581
rect -600 547 -432 581
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect 432 547 600 581
rect 690 547 858 581
rect 948 547 1116 581
rect 1206 547 1374 581
rect 1464 547 1632 581
rect 1722 547 1890 581
rect -1890 37 -1722 71
rect -1632 37 -1464 71
rect -1374 37 -1206 71
rect -1116 37 -948 71
rect -858 37 -690 71
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect 690 37 858 71
rect 948 37 1116 71
rect 1206 37 1374 71
rect 1464 37 1632 71
rect 1722 37 1890 71
rect -1890 -71 -1722 -37
rect -1632 -71 -1464 -37
rect -1374 -71 -1206 -37
rect -1116 -71 -948 -37
rect -858 -71 -690 -37
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect 690 -71 858 -37
rect 948 -71 1116 -37
rect 1206 -71 1374 -37
rect 1464 -71 1632 -37
rect 1722 -71 1890 -37
rect -1890 -581 -1722 -547
rect -1632 -581 -1464 -547
rect -1374 -581 -1206 -547
rect -1116 -581 -948 -547
rect -858 -581 -690 -547
rect -600 -581 -432 -547
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
rect 432 -581 600 -547
rect 690 -581 858 -547
rect 948 -581 1116 -547
rect 1206 -581 1374 -547
rect 1464 -581 1632 -547
rect 1722 -581 1890 -547
<< locali >>
rect -2066 587 -2032 683
rect 2032 587 2066 683
rect -1906 547 -1890 581
rect -1722 547 -1706 581
rect -1648 547 -1632 581
rect -1464 547 -1448 581
rect -1390 547 -1374 581
rect -1206 547 -1190 581
rect -1132 547 -1116 581
rect -948 547 -932 581
rect -874 547 -858 581
rect -690 547 -674 581
rect -616 547 -600 581
rect -432 547 -416 581
rect -358 547 -342 581
rect -174 547 -158 581
rect -100 547 -84 581
rect 84 547 100 581
rect 158 547 174 581
rect 342 547 358 581
rect 416 547 432 581
rect 600 547 616 581
rect 674 547 690 581
rect 858 547 874 581
rect 932 547 948 581
rect 1116 547 1132 581
rect 1190 547 1206 581
rect 1374 547 1390 581
rect 1448 547 1464 581
rect 1632 547 1648 581
rect 1706 547 1722 581
rect 1890 547 1906 581
rect -1952 497 -1918 513
rect -1952 105 -1918 121
rect -1694 497 -1660 513
rect -1694 105 -1660 121
rect -1436 497 -1402 513
rect -1436 105 -1402 121
rect -1178 497 -1144 513
rect -1178 105 -1144 121
rect -920 497 -886 513
rect -920 105 -886 121
rect -662 497 -628 513
rect -662 105 -628 121
rect -404 497 -370 513
rect -404 105 -370 121
rect -146 497 -112 513
rect -146 105 -112 121
rect 112 497 146 513
rect 112 105 146 121
rect 370 497 404 513
rect 370 105 404 121
rect 628 497 662 513
rect 628 105 662 121
rect 886 497 920 513
rect 886 105 920 121
rect 1144 497 1178 513
rect 1144 105 1178 121
rect 1402 497 1436 513
rect 1402 105 1436 121
rect 1660 497 1694 513
rect 1660 105 1694 121
rect 1918 497 1952 513
rect 1918 105 1952 121
rect -1906 37 -1890 71
rect -1722 37 -1706 71
rect -1648 37 -1632 71
rect -1464 37 -1448 71
rect -1390 37 -1374 71
rect -1206 37 -1190 71
rect -1132 37 -1116 71
rect -948 37 -932 71
rect -874 37 -858 71
rect -690 37 -674 71
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect 674 37 690 71
rect 858 37 874 71
rect 932 37 948 71
rect 1116 37 1132 71
rect 1190 37 1206 71
rect 1374 37 1390 71
rect 1448 37 1464 71
rect 1632 37 1648 71
rect 1706 37 1722 71
rect 1890 37 1906 71
rect -1906 -71 -1890 -37
rect -1722 -71 -1706 -37
rect -1648 -71 -1632 -37
rect -1464 -71 -1448 -37
rect -1390 -71 -1374 -37
rect -1206 -71 -1190 -37
rect -1132 -71 -1116 -37
rect -948 -71 -932 -37
rect -874 -71 -858 -37
rect -690 -71 -674 -37
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 416 -71 432 -37
rect 600 -71 616 -37
rect 674 -71 690 -37
rect 858 -71 874 -37
rect 932 -71 948 -37
rect 1116 -71 1132 -37
rect 1190 -71 1206 -37
rect 1374 -71 1390 -37
rect 1448 -71 1464 -37
rect 1632 -71 1648 -37
rect 1706 -71 1722 -37
rect 1890 -71 1906 -37
rect -1952 -121 -1918 -105
rect -1952 -513 -1918 -497
rect -1694 -121 -1660 -105
rect -1694 -513 -1660 -497
rect -1436 -121 -1402 -105
rect -1436 -513 -1402 -497
rect -1178 -121 -1144 -105
rect -1178 -513 -1144 -497
rect -920 -121 -886 -105
rect -920 -513 -886 -497
rect -662 -121 -628 -105
rect -662 -513 -628 -497
rect -404 -121 -370 -105
rect -404 -513 -370 -497
rect -146 -121 -112 -105
rect -146 -513 -112 -497
rect 112 -121 146 -105
rect 112 -513 146 -497
rect 370 -121 404 -105
rect 370 -513 404 -497
rect 628 -121 662 -105
rect 628 -513 662 -497
rect 886 -121 920 -105
rect 886 -513 920 -497
rect 1144 -121 1178 -105
rect 1144 -513 1178 -497
rect 1402 -121 1436 -105
rect 1402 -513 1436 -497
rect 1660 -121 1694 -105
rect 1660 -513 1694 -497
rect 1918 -121 1952 -105
rect 1918 -513 1952 -497
rect -1906 -581 -1890 -547
rect -1722 -581 -1706 -547
rect -1648 -581 -1632 -547
rect -1464 -581 -1448 -547
rect -1390 -581 -1374 -547
rect -1206 -581 -1190 -547
rect -1132 -581 -1116 -547
rect -948 -581 -932 -547
rect -874 -581 -858 -547
rect -690 -581 -674 -547
rect -616 -581 -600 -547
rect -432 -581 -416 -547
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 416 -581 432 -547
rect 600 -581 616 -547
rect 674 -581 690 -547
rect 858 -581 874 -547
rect 932 -581 948 -547
rect 1116 -581 1132 -547
rect 1190 -581 1206 -547
rect 1374 -581 1390 -547
rect 1448 -581 1464 -547
rect 1632 -581 1648 -547
rect 1706 -581 1722 -547
rect 1890 -581 1906 -547
rect -2066 -683 -1970 -649
rect 1970 -683 2066 -649
<< viali >>
rect -2032 649 2032 683
rect -1890 547 -1722 581
rect -1632 547 -1464 581
rect -1374 547 -1206 581
rect -1116 547 -948 581
rect -858 547 -690 581
rect -600 547 -432 581
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect 432 547 600 581
rect 690 547 858 581
rect 948 547 1116 581
rect 1206 547 1374 581
rect 1464 547 1632 581
rect 1722 547 1890 581
rect -1952 330 -1918 480
rect -1694 138 -1660 288
rect -1436 330 -1402 480
rect -1178 138 -1144 288
rect -920 330 -886 480
rect -662 138 -628 288
rect -404 330 -370 480
rect -146 138 -112 288
rect 112 330 146 480
rect 370 138 404 288
rect 628 330 662 480
rect 886 138 920 288
rect 1144 330 1178 480
rect 1402 138 1436 288
rect 1660 330 1694 480
rect 1918 138 1952 288
rect -1890 37 -1722 71
rect -1632 37 -1464 71
rect -1374 37 -1206 71
rect -1116 37 -948 71
rect -858 37 -690 71
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect 690 37 858 71
rect 948 37 1116 71
rect 1206 37 1374 71
rect 1464 37 1632 71
rect 1722 37 1890 71
rect -1890 -71 -1722 -37
rect -1632 -71 -1464 -37
rect -1374 -71 -1206 -37
rect -1116 -71 -948 -37
rect -858 -71 -690 -37
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect 690 -71 858 -37
rect 948 -71 1116 -37
rect 1206 -71 1374 -37
rect 1464 -71 1632 -37
rect 1722 -71 1890 -37
rect -2066 -587 -2032 -130
rect -1952 -288 -1918 -138
rect -1694 -480 -1660 -330
rect -1436 -288 -1402 -138
rect -1178 -480 -1144 -330
rect -920 -288 -886 -138
rect -662 -480 -628 -330
rect -404 -288 -370 -138
rect -146 -480 -112 -330
rect 112 -288 146 -138
rect 370 -480 404 -330
rect 628 -288 662 -138
rect 886 -480 920 -330
rect 1144 -288 1178 -138
rect 1402 -480 1436 -330
rect 1660 -288 1694 -138
rect 1918 -480 1952 -330
rect -1890 -581 -1722 -547
rect -1632 -581 -1464 -547
rect -1374 -581 -1206 -547
rect -1116 -581 -948 -547
rect -858 -581 -690 -547
rect -600 -581 -432 -547
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
rect 432 -581 600 -547
rect 690 -581 858 -547
rect 948 -581 1116 -547
rect 1206 -581 1374 -547
rect 1464 -581 1632 -547
rect 1722 -581 1890 -547
rect -2066 -649 -2032 -587
rect 2032 -587 2066 -130
rect 2032 -649 2066 -587
<< metal1 >>
rect -2044 683 2044 689
rect -2044 649 -2032 683
rect 2032 649 2044 683
rect -2044 643 2044 649
rect -1902 581 -1710 587
rect -1902 547 -1890 581
rect -1722 547 -1710 581
rect -1902 541 -1710 547
rect -1644 581 -1452 587
rect -1644 547 -1632 581
rect -1464 547 -1452 581
rect -1644 541 -1452 547
rect -1386 581 -1194 587
rect -1386 547 -1374 581
rect -1206 547 -1194 581
rect -1386 541 -1194 547
rect -1128 581 -936 587
rect -1128 547 -1116 581
rect -948 547 -936 581
rect -1128 541 -936 547
rect -870 581 -678 587
rect -870 547 -858 581
rect -690 547 -678 581
rect -870 541 -678 547
rect -612 581 -420 587
rect -612 547 -600 581
rect -432 547 -420 581
rect -612 541 -420 547
rect -354 581 -162 587
rect -354 547 -342 581
rect -174 547 -162 581
rect -354 541 -162 547
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect 162 581 354 587
rect 162 547 174 581
rect 342 547 354 581
rect 162 541 354 547
rect 420 581 612 587
rect 420 547 432 581
rect 600 547 612 581
rect 420 541 612 547
rect 678 581 870 587
rect 678 547 690 581
rect 858 547 870 581
rect 678 541 870 547
rect 936 581 1128 587
rect 936 547 948 581
rect 1116 547 1128 581
rect 936 541 1128 547
rect 1194 581 1386 587
rect 1194 547 1206 581
rect 1374 547 1386 581
rect 1194 541 1386 547
rect 1452 581 1644 587
rect 1452 547 1464 581
rect 1632 547 1644 581
rect 1452 541 1644 547
rect 1710 581 1902 587
rect 1710 547 1722 581
rect 1890 547 1902 581
rect 1710 541 1902 547
rect -1958 480 -1912 492
rect -1958 330 -1952 480
rect -1918 330 -1912 480
rect -1958 318 -1912 330
rect -1442 480 -1396 492
rect -1442 330 -1436 480
rect -1402 330 -1396 480
rect -1442 318 -1396 330
rect -926 480 -880 492
rect -926 330 -920 480
rect -886 330 -880 480
rect -926 318 -880 330
rect -410 480 -364 492
rect -410 330 -404 480
rect -370 330 -364 480
rect -410 318 -364 330
rect 106 480 152 492
rect 106 330 112 480
rect 146 330 152 480
rect 106 318 152 330
rect 622 480 668 492
rect 622 330 628 480
rect 662 330 668 480
rect 622 318 668 330
rect 1138 480 1184 492
rect 1138 330 1144 480
rect 1178 330 1184 480
rect 1138 318 1184 330
rect 1654 480 1700 492
rect 1654 330 1660 480
rect 1694 330 1700 480
rect 1654 318 1700 330
rect -1700 288 -1654 300
rect -1700 138 -1694 288
rect -1660 138 -1654 288
rect -1700 126 -1654 138
rect -1184 288 -1138 300
rect -1184 138 -1178 288
rect -1144 138 -1138 288
rect -1184 126 -1138 138
rect -668 288 -622 300
rect -668 138 -662 288
rect -628 138 -622 288
rect -668 126 -622 138
rect -152 288 -106 300
rect -152 138 -146 288
rect -112 138 -106 288
rect -152 126 -106 138
rect 364 288 410 300
rect 364 138 370 288
rect 404 138 410 288
rect 364 126 410 138
rect 880 288 926 300
rect 880 138 886 288
rect 920 138 926 288
rect 880 126 926 138
rect 1396 288 1442 300
rect 1396 138 1402 288
rect 1436 138 1442 288
rect 1396 126 1442 138
rect 1912 288 1958 300
rect 1912 138 1918 288
rect 1952 138 1958 288
rect 1912 126 1958 138
rect -1902 71 -1710 77
rect -1902 37 -1890 71
rect -1722 37 -1710 71
rect -1902 31 -1710 37
rect -1644 71 -1452 77
rect -1644 37 -1632 71
rect -1464 37 -1452 71
rect -1644 31 -1452 37
rect -1386 71 -1194 77
rect -1386 37 -1374 71
rect -1206 37 -1194 71
rect -1386 31 -1194 37
rect -1128 71 -936 77
rect -1128 37 -1116 71
rect -948 37 -936 71
rect -1128 31 -936 37
rect -870 71 -678 77
rect -870 37 -858 71
rect -690 37 -678 71
rect -870 31 -678 37
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect 678 71 870 77
rect 678 37 690 71
rect 858 37 870 71
rect 678 31 870 37
rect 936 71 1128 77
rect 936 37 948 71
rect 1116 37 1128 71
rect 936 31 1128 37
rect 1194 71 1386 77
rect 1194 37 1206 71
rect 1374 37 1386 71
rect 1194 31 1386 37
rect 1452 71 1644 77
rect 1452 37 1464 71
rect 1632 37 1644 71
rect 1452 31 1644 37
rect 1710 71 1902 77
rect 1710 37 1722 71
rect 1890 37 1902 71
rect 1710 31 1902 37
rect -1902 -37 -1710 -31
rect -1902 -71 -1890 -37
rect -1722 -71 -1710 -37
rect -1902 -77 -1710 -71
rect -1644 -37 -1452 -31
rect -1644 -71 -1632 -37
rect -1464 -71 -1452 -37
rect -1644 -77 -1452 -71
rect -1386 -37 -1194 -31
rect -1386 -71 -1374 -37
rect -1206 -71 -1194 -37
rect -1386 -77 -1194 -71
rect -1128 -37 -936 -31
rect -1128 -71 -1116 -37
rect -948 -71 -936 -37
rect -1128 -77 -936 -71
rect -870 -37 -678 -31
rect -870 -71 -858 -37
rect -690 -71 -678 -37
rect -870 -77 -678 -71
rect -612 -37 -420 -31
rect -612 -71 -600 -37
rect -432 -71 -420 -37
rect -612 -77 -420 -71
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect 420 -37 612 -31
rect 420 -71 432 -37
rect 600 -71 612 -37
rect 420 -77 612 -71
rect 678 -37 870 -31
rect 678 -71 690 -37
rect 858 -71 870 -37
rect 678 -77 870 -71
rect 936 -37 1128 -31
rect 936 -71 948 -37
rect 1116 -71 1128 -37
rect 936 -77 1128 -71
rect 1194 -37 1386 -31
rect 1194 -71 1206 -37
rect 1374 -71 1386 -37
rect 1194 -77 1386 -71
rect 1452 -37 1644 -31
rect 1452 -71 1464 -37
rect 1632 -71 1644 -37
rect 1452 -77 1644 -71
rect 1710 -37 1902 -31
rect 1710 -71 1722 -37
rect 1890 -71 1902 -37
rect 1710 -77 1902 -71
rect -2072 -130 -2026 -118
rect -2072 -649 -2066 -130
rect -2032 -649 -2026 -130
rect -1958 -138 -1912 -126
rect -1958 -288 -1952 -138
rect -1918 -288 -1912 -138
rect -1958 -300 -1912 -288
rect -1442 -138 -1396 -126
rect -1442 -288 -1436 -138
rect -1402 -288 -1396 -138
rect -1442 -300 -1396 -288
rect -926 -138 -880 -126
rect -926 -288 -920 -138
rect -886 -288 -880 -138
rect -926 -300 -880 -288
rect -410 -138 -364 -126
rect -410 -288 -404 -138
rect -370 -288 -364 -138
rect -410 -300 -364 -288
rect 106 -138 152 -126
rect 106 -288 112 -138
rect 146 -288 152 -138
rect 106 -300 152 -288
rect 622 -138 668 -126
rect 622 -288 628 -138
rect 662 -288 668 -138
rect 622 -300 668 -288
rect 1138 -138 1184 -126
rect 1138 -288 1144 -138
rect 1178 -288 1184 -138
rect 1138 -300 1184 -288
rect 1654 -138 1700 -126
rect 1654 -288 1660 -138
rect 1694 -288 1700 -138
rect 1654 -300 1700 -288
rect 2026 -130 2072 -118
rect -1700 -330 -1654 -318
rect -1700 -480 -1694 -330
rect -1660 -480 -1654 -330
rect -1700 -492 -1654 -480
rect -1184 -330 -1138 -318
rect -1184 -480 -1178 -330
rect -1144 -480 -1138 -330
rect -1184 -492 -1138 -480
rect -668 -330 -622 -318
rect -668 -480 -662 -330
rect -628 -480 -622 -330
rect -668 -492 -622 -480
rect -152 -330 -106 -318
rect -152 -480 -146 -330
rect -112 -480 -106 -330
rect -152 -492 -106 -480
rect 364 -330 410 -318
rect 364 -480 370 -330
rect 404 -480 410 -330
rect 364 -492 410 -480
rect 880 -330 926 -318
rect 880 -480 886 -330
rect 920 -480 926 -330
rect 880 -492 926 -480
rect 1396 -330 1442 -318
rect 1396 -480 1402 -330
rect 1436 -480 1442 -330
rect 1396 -492 1442 -480
rect 1912 -330 1958 -318
rect 1912 -480 1918 -330
rect 1952 -480 1958 -330
rect 1912 -492 1958 -480
rect -1902 -547 -1710 -541
rect -1902 -581 -1890 -547
rect -1722 -581 -1710 -547
rect -1902 -587 -1710 -581
rect -1644 -547 -1452 -541
rect -1644 -581 -1632 -547
rect -1464 -581 -1452 -547
rect -1644 -587 -1452 -581
rect -1386 -547 -1194 -541
rect -1386 -581 -1374 -547
rect -1206 -581 -1194 -547
rect -1386 -587 -1194 -581
rect -1128 -547 -936 -541
rect -1128 -581 -1116 -547
rect -948 -581 -936 -547
rect -1128 -587 -936 -581
rect -870 -547 -678 -541
rect -870 -581 -858 -547
rect -690 -581 -678 -547
rect -870 -587 -678 -581
rect -612 -547 -420 -541
rect -612 -581 -600 -547
rect -432 -581 -420 -547
rect -612 -587 -420 -581
rect -354 -547 -162 -541
rect -354 -581 -342 -547
rect -174 -581 -162 -547
rect -354 -587 -162 -581
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
rect 162 -547 354 -541
rect 162 -581 174 -547
rect 342 -581 354 -547
rect 162 -587 354 -581
rect 420 -547 612 -541
rect 420 -581 432 -547
rect 600 -581 612 -547
rect 420 -587 612 -581
rect 678 -547 870 -541
rect 678 -581 690 -547
rect 858 -581 870 -547
rect 678 -587 870 -581
rect 936 -547 1128 -541
rect 936 -581 948 -547
rect 1116 -581 1128 -547
rect 936 -587 1128 -581
rect 1194 -547 1386 -541
rect 1194 -581 1206 -547
rect 1374 -581 1386 -547
rect 1194 -587 1386 -581
rect 1452 -547 1644 -541
rect 1452 -581 1464 -547
rect 1632 -581 1644 -547
rect 1452 -587 1644 -581
rect 1710 -547 1902 -541
rect 1710 -581 1722 -547
rect 1890 -581 1902 -547
rect 1710 -587 1902 -581
rect -2072 -661 -2026 -649
rect 2026 -649 2032 -130
rect 2066 -649 2072 -130
rect 2026 -661 2072 -649
<< properties >>
string FIXED_BBOX -2049 -666 2049 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
