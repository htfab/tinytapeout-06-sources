magic
tech sky130A
magscale 1 2
timestamp 1710089296
<< viali >>
rect 3985 18921 4019 18955
rect 8493 18853 8527 18887
rect 9413 18785 9447 18819
rect 15577 18785 15611 18819
rect 16221 18785 16255 18819
rect 18153 18785 18187 18819
rect 857 18717 891 18751
rect 9137 18717 9171 18751
rect 9321 18717 9355 18751
rect 8677 18649 8711 18683
rect 9781 18581 9815 18615
rect 10793 18241 10827 18275
rect 6377 18173 6411 18207
rect 6653 18105 6687 18139
rect 10517 18105 10551 18139
rect 8125 18037 8159 18071
rect 9045 18037 9079 18071
rect 10057 17833 10091 17867
rect 11161 17833 11195 17867
rect 6713 17765 6747 17799
rect 6929 17765 6963 17799
rect 7481 17765 7515 17799
rect 11529 17765 11563 17799
rect 5641 17697 5675 17731
rect 6469 17697 6503 17731
rect 9873 17697 9907 17731
rect 10977 17697 11011 17731
rect 3617 17629 3651 17663
rect 3893 17629 3927 17663
rect 7205 17629 7239 17663
rect 11253 17629 11287 17663
rect 5825 17493 5859 17527
rect 6561 17493 6595 17527
rect 6745 17493 6779 17527
rect 8953 17493 8987 17527
rect 13001 17493 13035 17527
rect 4445 17289 4479 17323
rect 4813 17289 4847 17323
rect 6101 17289 6135 17323
rect 7297 17289 7331 17323
rect 11437 17289 11471 17323
rect 4997 17221 5031 17255
rect 6193 17221 6227 17255
rect 7665 17221 7699 17255
rect 6469 17153 6503 17187
rect 11989 17153 12023 17187
rect 4629 17085 4663 17119
rect 4905 17085 4939 17119
rect 5273 17085 5307 17119
rect 6285 17085 6319 17119
rect 6377 17085 6411 17119
rect 6561 17085 6595 17119
rect 6653 17085 6687 17119
rect 6837 17085 6871 17119
rect 6929 17085 6963 17119
rect 7021 17085 7055 17119
rect 7389 17085 7423 17119
rect 8769 17085 8803 17119
rect 9045 17085 9079 17119
rect 11897 17085 11931 17119
rect 4997 17017 5031 17051
rect 6009 17017 6043 17051
rect 7665 17017 7699 17051
rect 9321 17017 9355 17051
rect 5181 16949 5215 16983
rect 7481 16949 7515 16983
rect 8953 16949 8987 16983
rect 10793 16949 10827 16983
rect 11805 16949 11839 16983
rect 7113 16745 7147 16779
rect 8585 16745 8619 16779
rect 9045 16745 9079 16779
rect 7481 16677 7515 16711
rect 8953 16677 8987 16711
rect 7251 16643 7285 16677
rect 3709 16609 3743 16643
rect 5273 16609 5307 16643
rect 6653 16609 6687 16643
rect 6745 16609 6779 16643
rect 6837 16609 6871 16643
rect 7021 16609 7055 16643
rect 18797 16609 18831 16643
rect 18981 16609 19015 16643
rect 9137 16541 9171 16575
rect 3525 16405 3559 16439
rect 5549 16405 5583 16439
rect 6377 16405 6411 16439
rect 7297 16405 7331 16439
rect 7297 16201 7331 16235
rect 4997 16133 5031 16167
rect 12449 16133 12483 16167
rect 3249 16065 3283 16099
rect 9045 16065 9079 16099
rect 9873 16065 9907 16099
rect 11805 16065 11839 16099
rect 7205 15997 7239 16031
rect 7849 15997 7883 16031
rect 9597 15997 9631 16031
rect 11989 15997 12023 16031
rect 12725 15997 12759 16031
rect 18981 15997 19015 16031
rect 3525 15929 3559 15963
rect 10149 15929 10183 15963
rect 6561 15861 6595 15895
rect 8401 15861 8435 15895
rect 8769 15861 8803 15895
rect 8861 15861 8895 15895
rect 9781 15861 9815 15895
rect 11621 15861 11655 15895
rect 12081 15861 12115 15895
rect 12541 15861 12575 15895
rect 18797 15861 18831 15895
rect 5917 15657 5951 15691
rect 9965 15657 9999 15691
rect 10425 15657 10459 15691
rect 13461 15657 13495 15691
rect 3785 15589 3819 15623
rect 3985 15589 4019 15623
rect 6377 15589 6411 15623
rect 8217 15589 8251 15623
rect 11989 15589 12023 15623
rect 2881 15521 2915 15555
rect 4353 15521 4387 15555
rect 5457 15521 5491 15555
rect 5549 15521 5583 15555
rect 5825 15521 5859 15555
rect 6009 15521 6043 15555
rect 6101 15521 6135 15555
rect 7941 15521 7975 15555
rect 10333 15521 10367 15555
rect 11713 15521 11747 15555
rect 18613 15521 18647 15555
rect 5273 15453 5307 15487
rect 5365 15453 5399 15487
rect 9689 15453 9723 15487
rect 10517 15453 10551 15487
rect 17509 15453 17543 15487
rect 18521 15453 18555 15487
rect 3617 15385 3651 15419
rect 2329 15317 2363 15351
rect 3801 15317 3835 15351
rect 4261 15317 4295 15351
rect 5089 15317 5123 15351
rect 7849 15317 7883 15351
rect 3893 15113 3927 15147
rect 4629 15113 4663 15147
rect 6837 15113 6871 15147
rect 7021 15113 7055 15147
rect 8217 15113 8251 15147
rect 8769 15045 8803 15079
rect 18337 15045 18371 15079
rect 2881 14977 2915 15011
rect 3525 14977 3559 15011
rect 4997 14977 5031 15011
rect 6745 14977 6779 15011
rect 16865 14977 16899 15011
rect 857 14909 891 14943
rect 3249 14909 3283 14943
rect 3341 14909 3375 14943
rect 4077 14909 4111 14943
rect 4169 14909 4203 14943
rect 4261 14909 4295 14943
rect 4353 14909 4387 14943
rect 4813 14909 4847 14943
rect 8033 14909 8067 14943
rect 9137 14909 9171 14943
rect 11345 14909 11379 14943
rect 11621 14909 11655 14943
rect 18337 14909 18371 14943
rect 1133 14841 1167 14875
rect 5273 14841 5307 14875
rect 7205 14841 7239 14875
rect 8493 14841 8527 14875
rect 9413 14841 9447 14875
rect 11897 14841 11931 14875
rect 18797 14841 18831 14875
rect 18981 14841 19015 14875
rect 3525 14773 3559 14807
rect 7005 14773 7039 14807
rect 10885 14773 10919 14807
rect 11529 14773 11563 14807
rect 13369 14773 13403 14807
rect 1409 14569 1443 14603
rect 2145 14569 2179 14603
rect 4629 14569 4663 14603
rect 4813 14569 4847 14603
rect 6193 14569 6227 14603
rect 9045 14569 9079 14603
rect 9597 14569 9631 14603
rect 11713 14569 11747 14603
rect 14933 14569 14967 14603
rect 4445 14501 4479 14535
rect 5825 14501 5859 14535
rect 6285 14501 6319 14535
rect 15025 14501 15059 14535
rect 1593 14433 1627 14467
rect 1869 14433 1903 14467
rect 1961 14433 1995 14467
rect 2237 14433 2271 14467
rect 2329 14433 2363 14467
rect 4537 14433 4571 14467
rect 6561 14433 6595 14467
rect 7757 14433 7791 14467
rect 9781 14433 9815 14467
rect 12081 14433 12115 14467
rect 12173 14433 12207 14467
rect 14381 14433 14415 14467
rect 15117 14433 15151 14467
rect 15577 14433 15611 14467
rect 16313 14433 16347 14467
rect 16497 14433 16531 14467
rect 16865 14433 16899 14467
rect 18337 14433 18371 14467
rect 18981 14433 19015 14467
rect 1777 14365 1811 14399
rect 2605 14365 2639 14399
rect 5917 14365 5951 14399
rect 12265 14365 12299 14399
rect 14565 14365 14599 14399
rect 15761 14365 15795 14399
rect 16129 14365 16163 14399
rect 16957 14365 16991 14399
rect 1961 14297 1995 14331
rect 4077 14297 4111 14331
rect 4261 14297 4295 14331
rect 18245 14297 18279 14331
rect 6009 14229 6043 14263
rect 6469 14229 6503 14263
rect 15393 14229 15427 14263
rect 16681 14229 16715 14263
rect 18705 14229 18739 14263
rect 2789 14025 2823 14059
rect 4905 14025 4939 14059
rect 6377 14025 6411 14059
rect 9413 14025 9447 14059
rect 14381 14025 14415 14059
rect 18889 14025 18923 14059
rect 3249 13957 3283 13991
rect 6929 13957 6963 13991
rect 10793 13957 10827 13991
rect 15117 13957 15151 13991
rect 9965 13889 9999 13923
rect 14657 13889 14691 13923
rect 16773 13889 16807 13923
rect 17049 13889 17083 13923
rect 2605 13821 2639 13855
rect 2789 13821 2823 13855
rect 3433 13821 3467 13855
rect 3617 13821 3651 13855
rect 6193 13821 6227 13855
rect 7205 13821 7239 13855
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 10241 13821 10275 13855
rect 10517 13821 10551 13855
rect 10609 13821 10643 13855
rect 11253 13821 11287 13855
rect 12449 13821 12483 13855
rect 14565 13821 14599 13855
rect 15301 13821 15335 13855
rect 16865 13821 16899 13855
rect 17233 13821 17267 13855
rect 18521 13821 18555 13855
rect 19073 13821 19107 13855
rect 6561 13753 6595 13787
rect 6653 13753 6687 13787
rect 10425 13753 10459 13787
rect 11069 13753 11103 13787
rect 12265 13753 12299 13787
rect 15117 13753 15151 13787
rect 6745 13685 6779 13719
rect 7021 13685 7055 13719
rect 10885 13685 10919 13719
rect 12081 13685 12115 13719
rect 5473 13481 5507 13515
rect 5993 13481 6027 13515
rect 8677 13481 8711 13515
rect 13553 13481 13587 13515
rect 13737 13481 13771 13515
rect 17969 13481 18003 13515
rect 5273 13413 5307 13447
rect 6193 13413 6227 13447
rect 6837 13413 6871 13447
rect 9137 13413 9171 13447
rect 12081 13413 12115 13447
rect 14289 13413 14323 13447
rect 1961 13345 1995 13379
rect 5181 13345 5215 13379
rect 6561 13345 6595 13379
rect 8493 13345 8527 13379
rect 8677 13345 8711 13379
rect 8850 13345 8884 13379
rect 8954 13345 8988 13379
rect 9229 13345 9263 13379
rect 9345 13345 9379 13379
rect 9597 13345 9631 13379
rect 9781 13345 9815 13379
rect 10149 13345 10183 13379
rect 11161 13345 11195 13379
rect 11254 13345 11288 13379
rect 11437 13345 11471 13379
rect 11529 13345 11563 13379
rect 11667 13345 11701 13379
rect 11897 13345 11931 13379
rect 12173 13345 12207 13379
rect 12265 13345 12299 13379
rect 12909 13345 12943 13379
rect 13001 13345 13035 13379
rect 13093 13345 13127 13379
rect 13211 13345 13245 13379
rect 13369 13345 13403 13379
rect 14473 13345 14507 13379
rect 15025 13345 15059 13379
rect 15577 13345 15611 13379
rect 15669 13345 15703 13379
rect 16129 13345 16163 13379
rect 17601 13345 17635 13379
rect 18245 13345 18279 13379
rect 1685 13277 1719 13311
rect 4905 13277 4939 13311
rect 10057 13277 10091 13311
rect 10793 13277 10827 13311
rect 13829 13277 13863 13311
rect 1869 13209 1903 13243
rect 5641 13209 5675 13243
rect 14289 13209 14323 13243
rect 17601 13209 17635 13243
rect 1777 13141 1811 13175
rect 4261 13141 4295 13175
rect 4997 13141 5031 13175
rect 5457 13141 5491 13175
rect 5825 13141 5859 13175
rect 6009 13141 6043 13175
rect 8309 13141 8343 13175
rect 9505 13141 9539 13175
rect 11805 13141 11839 13175
rect 12449 13141 12483 13175
rect 12725 13141 12759 13175
rect 14565 13141 14599 13175
rect 18613 13141 18647 13175
rect 2605 12937 2639 12971
rect 2881 12937 2915 12971
rect 6193 12937 6227 12971
rect 7205 12937 7239 12971
rect 10241 12937 10275 12971
rect 11621 12937 11655 12971
rect 12541 12937 12575 12971
rect 12633 12937 12667 12971
rect 11161 12869 11195 12903
rect 1133 12801 1167 12835
rect 4353 12801 4387 12835
rect 4629 12801 4663 12835
rect 6101 12801 6135 12835
rect 6653 12801 6687 12835
rect 6837 12801 6871 12835
rect 7665 12801 7699 12835
rect 7849 12801 7883 12835
rect 10057 12801 10091 12835
rect 11437 12801 11471 12835
rect 14080 12801 14114 12835
rect 14197 12801 14231 12835
rect 14565 12801 14599 12835
rect 15025 12801 15059 12835
rect 16221 12801 16255 12835
rect 17785 12801 17819 12835
rect 19073 12801 19107 12835
rect 857 12733 891 12767
rect 3525 12733 3559 12767
rect 3617 12733 3651 12767
rect 3709 12733 3743 12767
rect 3893 12733 3927 12767
rect 8585 12733 8619 12767
rect 8678 12733 8712 12767
rect 9050 12733 9084 12767
rect 9321 12733 9355 12767
rect 9505 12733 9539 12767
rect 9921 12733 9955 12767
rect 10609 12733 10643 12767
rect 10885 12733 10919 12767
rect 10977 12733 11011 12767
rect 11345 12733 11379 12767
rect 11621 12733 11655 12767
rect 12725 12733 12759 12767
rect 12817 12733 12851 12767
rect 13001 12733 13035 12767
rect 15117 12733 15151 12767
rect 16313 12733 16347 12767
rect 17877 12733 17911 12767
rect 18705 12733 18739 12767
rect 2697 12665 2731 12699
rect 2913 12665 2947 12699
rect 7573 12665 7607 12699
rect 8861 12665 8895 12699
rect 8953 12665 8987 12699
rect 10793 12665 10827 12699
rect 13553 12665 13587 12699
rect 13737 12665 13771 12699
rect 3065 12597 3099 12631
rect 3249 12597 3283 12631
rect 6561 12597 6595 12631
rect 9229 12597 9263 12631
rect 11805 12597 11839 12631
rect 12265 12597 12299 12631
rect 13921 12597 13955 12631
rect 14289 12597 14323 12631
rect 18705 12597 18739 12631
rect 4905 12393 4939 12427
rect 8401 12393 8435 12427
rect 11805 12393 11839 12427
rect 11973 12393 12007 12427
rect 13185 12393 13219 12427
rect 13553 12393 13587 12427
rect 1869 12325 1903 12359
rect 2492 12325 2526 12359
rect 2697 12325 2731 12359
rect 3433 12325 3467 12359
rect 7389 12325 7423 12359
rect 9045 12325 9079 12359
rect 12173 12325 12207 12359
rect 13461 12325 13495 12359
rect 1777 12257 1811 12291
rect 2053 12257 2087 12291
rect 2789 12257 2823 12291
rect 2973 12257 3007 12291
rect 6469 12257 6503 12291
rect 7205 12257 7239 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 7849 12257 7883 12291
rect 8033 12257 8067 12291
rect 8125 12257 8159 12291
rect 8217 12257 8251 12291
rect 9505 12257 9539 12291
rect 9689 12257 9723 12291
rect 10057 12257 10091 12291
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 12449 12257 12483 12291
rect 13001 12257 13035 12291
rect 15485 12257 15519 12291
rect 16405 12257 16439 12291
rect 17877 12257 17911 12291
rect 2881 12189 2915 12223
rect 3157 12189 3191 12223
rect 9965 12189 9999 12223
rect 12725 12189 12759 12223
rect 12817 12189 12851 12223
rect 12909 12189 12943 12223
rect 13344 12189 13378 12223
rect 13829 12189 13863 12223
rect 14381 12189 14415 12223
rect 15393 12189 15427 12223
rect 16497 12189 16531 12223
rect 2053 12121 2087 12155
rect 11437 12121 11471 12155
rect 12265 12121 12299 12155
rect 17785 12121 17819 12155
rect 2329 12053 2363 12087
rect 2513 12053 2547 12087
rect 6285 12053 6319 12087
rect 7757 12053 7791 12087
rect 11989 12053 12023 12087
rect 12541 12053 12575 12087
rect 16221 12053 16255 12087
rect 4721 11849 4755 11883
rect 7573 11849 7607 11883
rect 10057 11849 10091 11883
rect 1501 11781 1535 11815
rect 2973 11781 3007 11815
rect 5825 11713 5859 11747
rect 6101 11713 6135 11747
rect 9413 11713 9447 11747
rect 9781 11713 9815 11747
rect 14289 11713 14323 11747
rect 16957 11713 16991 11747
rect 1501 11645 1535 11679
rect 1685 11645 1719 11679
rect 1777 11645 1811 11679
rect 2697 11645 2731 11679
rect 4445 11645 4479 11679
rect 4905 11645 4939 11679
rect 5181 11645 5215 11679
rect 8677 11645 8711 11679
rect 9321 11645 9355 11679
rect 9689 11645 9723 11679
rect 11069 11645 11103 11679
rect 11253 11645 11287 11679
rect 11621 11645 11655 11679
rect 11805 11645 11839 11679
rect 14197 11645 14231 11679
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 17049 11645 17083 11679
rect 17325 11645 17359 11679
rect 19073 11645 19107 11679
rect 2789 11577 2823 11611
rect 2973 11577 3007 11611
rect 8493 11577 8527 11611
rect 12265 11577 12299 11611
rect 17141 11577 17175 11611
rect 4353 11509 4387 11543
rect 4997 11509 5031 11543
rect 8861 11509 8895 11543
rect 18889 11509 18923 11543
rect 4905 11305 4939 11339
rect 5273 11305 5307 11339
rect 6469 11305 6503 11339
rect 6929 11305 6963 11339
rect 8309 11305 8343 11339
rect 6837 11237 6871 11271
rect 8769 11237 8803 11271
rect 10333 11237 10367 11271
rect 10425 11237 10459 11271
rect 13369 11237 13403 11271
rect 13829 11237 13863 11271
rect 14289 11237 14323 11271
rect 15117 11237 15151 11271
rect 18153 11237 18187 11271
rect 18889 11237 18923 11271
rect 857 11169 891 11203
rect 2881 11169 2915 11203
rect 5365 11169 5399 11203
rect 8125 11169 8159 11203
rect 8217 11169 8251 11203
rect 8493 11169 8527 11203
rect 9413 11169 9447 11203
rect 9781 11169 9815 11203
rect 9873 11169 9907 11203
rect 10057 11169 10091 11203
rect 10215 11169 10249 11203
rect 10517 11169 10551 11203
rect 10977 11169 11011 11203
rect 11253 11169 11287 11203
rect 11437 11169 11471 11203
rect 11805 11169 11839 11203
rect 12725 11169 12759 11203
rect 13001 11169 13035 11203
rect 14013 11169 14047 11203
rect 14197 11169 14231 11203
rect 14381 11169 14415 11203
rect 15393 11169 15427 11203
rect 16497 11169 16531 11203
rect 17785 11169 17819 11203
rect 1133 11101 1167 11135
rect 3157 11101 3191 11135
rect 5549 11101 5583 11135
rect 7021 11101 7055 11135
rect 9229 11101 9263 11135
rect 11069 11101 11103 11135
rect 11713 11101 11747 11135
rect 12449 11101 12483 11135
rect 13277 11101 13311 11135
rect 14933 11101 14967 11135
rect 15025 11101 15059 11135
rect 4629 11033 4663 11067
rect 8033 11033 8067 11067
rect 8677 11033 8711 11067
rect 10701 11033 10735 11067
rect 12541 11033 12575 11067
rect 12909 11033 12943 11067
rect 13093 11033 13127 11067
rect 13829 11033 13863 11067
rect 14565 11033 14599 11067
rect 17785 11033 17819 11067
rect 2605 10965 2639 10999
rect 14749 10965 14783 10999
rect 1317 10761 1351 10795
rect 3249 10761 3283 10795
rect 6009 10761 6043 10795
rect 10885 10761 10919 10795
rect 10977 10761 11011 10795
rect 3341 10693 3375 10727
rect 10793 10693 10827 10727
rect 13553 10693 13587 10727
rect 14289 10693 14323 10727
rect 2789 10625 2823 10659
rect 4261 10625 4295 10659
rect 8401 10625 8435 10659
rect 10333 10625 10367 10659
rect 13829 10625 13863 10659
rect 15853 10625 15887 10659
rect 16405 10625 16439 10659
rect 17877 10625 17911 10659
rect 1501 10557 1535 10591
rect 1685 10557 1719 10591
rect 1777 10557 1811 10591
rect 2237 10557 2271 10591
rect 3249 10557 3283 10591
rect 8861 10557 8895 10591
rect 9045 10557 9079 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 9689 10557 9723 10591
rect 9965 10557 9999 10591
rect 10149 10557 10183 10591
rect 10517 10557 10551 10591
rect 13737 10557 13771 10591
rect 14841 10557 14875 10591
rect 15209 10557 15243 10591
rect 15485 10557 15519 10591
rect 16129 10557 16163 10591
rect 16313 10557 16347 10591
rect 17969 10557 18003 10591
rect 18245 10557 18279 10591
rect 18889 10557 18923 10591
rect 3525 10489 3559 10523
rect 4537 10489 4571 10523
rect 9827 10489 9861 10523
rect 10057 10489 10091 10523
rect 14289 10489 14323 10523
rect 15577 10489 15611 10523
rect 15945 10489 15979 10523
rect 18337 10489 18371 10523
rect 10609 10421 10643 10455
rect 11253 10421 11287 10455
rect 18061 10421 18095 10455
rect 18705 10421 18739 10455
rect 3065 10217 3099 10251
rect 12173 10217 12207 10251
rect 12633 10217 12667 10251
rect 12817 10217 12851 10251
rect 14289 10217 14323 10251
rect 15393 10217 15427 10251
rect 2789 10149 2823 10183
rect 7205 10149 7239 10183
rect 9137 10149 9171 10183
rect 2973 10081 3007 10115
rect 3157 10081 3191 10115
rect 3341 10081 3375 10115
rect 3525 10081 3559 10115
rect 6653 10081 6687 10115
rect 9045 10081 9079 10115
rect 9321 10081 9355 10115
rect 9597 10081 9631 10115
rect 10149 10081 10183 10115
rect 10333 10081 10367 10115
rect 10425 10081 10459 10115
rect 10517 10081 10551 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 12357 10081 12391 10115
rect 13737 10081 13771 10115
rect 14381 10081 14415 10115
rect 15025 10081 15059 10115
rect 15209 10081 15243 10115
rect 15577 10081 15611 10115
rect 15669 10081 15703 10115
rect 15853 10081 15887 10115
rect 16497 10081 16531 10115
rect 16773 10081 16807 10115
rect 17141 10081 17175 10115
rect 17417 10081 17451 10115
rect 18521 10081 18555 10115
rect 9689 10013 9723 10047
rect 12541 10013 12575 10047
rect 14013 10013 14047 10047
rect 14498 10013 14532 10047
rect 16313 10013 16347 10047
rect 17325 10013 17359 10047
rect 18429 10013 18463 10047
rect 3709 9945 3743 9979
rect 9965 9945 9999 9979
rect 10701 9945 10735 9979
rect 13185 9945 13219 9979
rect 13461 9945 13495 9979
rect 16129 9945 16163 9979
rect 6469 9877 6503 9911
rect 8493 9877 8527 9911
rect 9505 9877 9539 9911
rect 9597 9877 9631 9911
rect 11069 9877 11103 9911
rect 11345 9877 11379 9911
rect 12817 9877 12851 9911
rect 13277 9877 13311 9911
rect 14657 9877 14691 9911
rect 15117 9877 15151 9911
rect 15761 9877 15795 9911
rect 16313 9877 16347 9911
rect 16405 9877 16439 9911
rect 16865 9877 16899 9911
rect 8401 9673 8435 9707
rect 10149 9673 10183 9707
rect 11529 9673 11563 9707
rect 12449 9673 12483 9707
rect 18245 9673 18279 9707
rect 18705 9673 18739 9707
rect 3249 9605 3283 9639
rect 10885 9605 10919 9639
rect 12357 9605 12391 9639
rect 17693 9605 17727 9639
rect 6009 9537 6043 9571
rect 6285 9537 6319 9571
rect 7757 9537 7791 9571
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 12541 9537 12575 9571
rect 15761 9537 15795 9571
rect 16037 9537 16071 9571
rect 19073 9537 19107 9571
rect 2421 9469 2455 9503
rect 2605 9469 2639 9503
rect 9505 9469 9539 9503
rect 9598 9469 9632 9503
rect 9781 9469 9815 9503
rect 10011 9469 10045 9503
rect 10241 9469 10275 9503
rect 10389 9469 10423 9503
rect 10517 9469 10551 9503
rect 10747 9469 10781 9503
rect 10977 9469 11011 9503
rect 11069 9469 11103 9503
rect 11253 9469 11287 9503
rect 11345 9469 11379 9503
rect 11713 9469 11747 9503
rect 11806 9469 11840 9503
rect 12081 9469 12115 9503
rect 12219 9469 12253 9503
rect 12449 9469 12483 9503
rect 14197 9469 14231 9503
rect 14473 9469 14507 9503
rect 14657 9469 14691 9503
rect 14933 9469 14967 9503
rect 15126 9469 15160 9503
rect 15945 9469 15979 9503
rect 17509 9469 17543 9503
rect 17601 9469 17635 9503
rect 17877 9469 17911 9503
rect 17969 9469 18003 9503
rect 18245 9469 18279 9503
rect 18429 9469 18463 9503
rect 18889 9469 18923 9503
rect 2789 9401 2823 9435
rect 3433 9401 3467 9435
rect 9873 9401 9907 9435
rect 10609 9401 10643 9435
rect 11989 9401 12023 9435
rect 8769 9333 8803 9367
rect 12817 9333 12851 9367
rect 18153 9333 18187 9367
rect 2697 9129 2731 9163
rect 4353 9129 4387 9163
rect 4813 9129 4847 9163
rect 5549 9129 5583 9163
rect 7573 9129 7607 9163
rect 8677 9129 8711 9163
rect 10333 9129 10367 9163
rect 11345 9129 11379 9163
rect 11805 9129 11839 9163
rect 15761 9129 15795 9163
rect 4537 9061 4571 9095
rect 6101 9061 6135 9095
rect 8309 9061 8343 9095
rect 9965 9061 9999 9095
rect 10977 9061 11011 9095
rect 11177 9061 11211 9095
rect 11437 9061 11471 9095
rect 11637 9061 11671 9095
rect 15577 9061 15611 9095
rect 16313 9061 16347 9095
rect 2881 8993 2915 9027
rect 3801 8993 3835 9027
rect 4077 8993 4111 9027
rect 4629 8993 4663 9027
rect 4905 8993 4939 9027
rect 5365 8993 5399 9027
rect 9689 8993 9723 9027
rect 9847 8993 9881 9027
rect 10057 8993 10091 9027
rect 10149 8993 10183 9027
rect 14105 8993 14139 9027
rect 14289 8993 14323 9027
rect 14381 8993 14415 9027
rect 14565 8993 14599 9027
rect 14933 8993 14967 9027
rect 15669 8993 15703 9027
rect 15853 8993 15887 9027
rect 16589 8993 16623 9027
rect 17049 8993 17083 9027
rect 17417 8993 17451 9027
rect 18613 8993 18647 9027
rect 857 8925 891 8959
rect 1133 8925 1167 8959
rect 3065 8925 3099 8959
rect 3525 8925 3559 8959
rect 5825 8925 5859 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 13553 8925 13587 8959
rect 14013 8925 14047 8959
rect 14841 8925 14875 8959
rect 17509 8925 17543 8959
rect 18521 8925 18555 8959
rect 3709 8857 3743 8891
rect 4629 8857 4663 8891
rect 13829 8857 13863 8891
rect 2605 8789 2639 8823
rect 3617 8789 3651 8823
rect 4353 8789 4387 8823
rect 11161 8789 11195 8823
rect 11621 8789 11655 8823
rect 14197 8789 14231 8823
rect 1501 8585 1535 8619
rect 3512 8585 3546 8619
rect 5733 8585 5767 8619
rect 8217 8585 8251 8619
rect 9505 8585 9539 8619
rect 12081 8585 12115 8619
rect 1593 8517 1627 8551
rect 2053 8517 2087 8551
rect 4997 8517 5031 8551
rect 13369 8517 13403 8551
rect 18429 8517 18463 8551
rect 3249 8449 3283 8483
rect 6193 8449 6227 8483
rect 6377 8449 6411 8483
rect 7665 8449 7699 8483
rect 8861 8449 8895 8483
rect 12173 8449 12207 8483
rect 14841 8449 14875 8483
rect 15393 8449 15427 8483
rect 16957 8449 16991 8483
rect 19073 8449 19107 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 1777 8381 1811 8415
rect 2053 8381 2087 8415
rect 6101 8381 6135 8415
rect 7849 8381 7883 8415
rect 9137 8381 9171 8415
rect 11437 8381 11471 8415
rect 11529 8381 11563 8415
rect 11713 8381 11747 8415
rect 11805 8381 11839 8415
rect 12357 8381 12391 8415
rect 12633 8381 12667 8415
rect 12817 8381 12851 8415
rect 13185 8381 13219 8415
rect 13737 8381 13771 8415
rect 13921 8381 13955 8415
rect 14197 8381 14231 8415
rect 14473 8381 14507 8415
rect 15209 8381 15243 8415
rect 15761 8381 15795 8415
rect 16865 8381 16899 8415
rect 18061 8381 18095 8415
rect 18889 8381 18923 8415
rect 1869 8313 1903 8347
rect 7757 8313 7791 8347
rect 11989 8313 12023 8347
rect 12081 8313 12115 8347
rect 14381 8313 14415 8347
rect 9045 8245 9079 8279
rect 12541 8245 12575 8279
rect 12909 8245 12943 8279
rect 18705 8245 18739 8279
rect 1869 8041 1903 8075
rect 7573 8041 7607 8075
rect 8401 8041 8435 8075
rect 9045 8041 9079 8075
rect 1685 7973 1719 8007
rect 8125 7973 8159 8007
rect 8677 7973 8711 8007
rect 8769 7973 8803 8007
rect 1961 7905 1995 7939
rect 5457 7905 5491 7939
rect 5825 7905 5859 7939
rect 7849 7905 7883 7939
rect 8033 7905 8067 7939
rect 8241 7905 8275 7939
rect 8493 7905 8527 7939
rect 8861 7905 8895 7939
rect 11713 7905 11747 7939
rect 11805 7905 11839 7939
rect 12173 7905 12207 7939
rect 12265 7905 12299 7939
rect 12633 7905 12667 7939
rect 13185 7905 13219 7939
rect 13645 7905 13679 7939
rect 14197 7905 14231 7939
rect 15117 7905 15151 7939
rect 15393 7905 15427 7939
rect 15945 7905 15979 7939
rect 16313 7905 16347 7939
rect 16405 7905 16439 7939
rect 16589 7905 16623 7939
rect 17693 7905 17727 7939
rect 18245 7905 18279 7939
rect 18521 7905 18555 7939
rect 18797 7905 18831 7939
rect 18981 7905 19015 7939
rect 6101 7837 6135 7871
rect 12725 7837 12759 7871
rect 12817 7837 12851 7871
rect 12909 7837 12943 7871
rect 14289 7837 14323 7871
rect 18613 7837 18647 7871
rect 5641 7769 5675 7803
rect 14565 7769 14599 7803
rect 15025 7769 15059 7803
rect 17877 7769 17911 7803
rect 1685 7701 1719 7735
rect 11253 7701 11287 7735
rect 13093 7701 13127 7735
rect 16129 7701 16163 7735
rect 2605 7497 2639 7531
rect 6193 7497 6227 7531
rect 8953 7497 8987 7531
rect 11897 7497 11931 7531
rect 6745 7429 6779 7463
rect 13737 7429 13771 7463
rect 857 7361 891 7395
rect 7297 7361 7331 7395
rect 9873 7361 9907 7395
rect 10333 7361 10367 7395
rect 13277 7361 13311 7395
rect 15393 7361 15427 7395
rect 17969 7361 18003 7395
rect 18705 7361 18739 7395
rect 19073 7361 19107 7395
rect 3985 7293 4019 7327
rect 4261 7293 4295 7327
rect 7113 7293 7147 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 9965 7293 9999 7327
rect 10149 7293 10183 7327
rect 10793 7293 10827 7327
rect 11437 7293 11471 7327
rect 11713 7293 11747 7327
rect 12449 7293 12483 7327
rect 12633 7293 12667 7327
rect 13185 7293 13219 7327
rect 13553 7293 13587 7327
rect 14289 7293 14323 7327
rect 15117 7293 15151 7327
rect 15761 7293 15795 7327
rect 16865 7293 16899 7327
rect 16957 7293 16991 7327
rect 18061 7293 18095 7327
rect 18889 7293 18923 7327
rect 1133 7225 1167 7259
rect 4905 7225 4939 7259
rect 9689 7225 9723 7259
rect 10885 7225 10919 7259
rect 12081 7225 12115 7259
rect 13829 7225 13863 7259
rect 3801 7157 3835 7191
rect 4169 7157 4203 7191
rect 7205 7157 7239 7191
rect 9965 7157 9999 7191
rect 10701 7157 10735 7191
rect 11529 7157 11563 7191
rect 10241 6953 10275 6987
rect 11621 6953 11655 6987
rect 3601 6885 3635 6919
rect 3801 6885 3835 6919
rect 10057 6885 10091 6919
rect 1685 6817 1719 6851
rect 1869 6817 1903 6851
rect 2973 6817 3007 6851
rect 3249 6817 3283 6851
rect 3893 6817 3927 6851
rect 4077 6817 4111 6851
rect 7941 6817 7975 6851
rect 10333 6817 10367 6851
rect 11713 6817 11747 6851
rect 11897 6817 11931 6851
rect 12357 6817 12391 6851
rect 12541 6817 12575 6851
rect 13277 6817 13311 6851
rect 14197 6817 14231 6851
rect 15853 6817 15887 6851
rect 16405 6817 16439 6851
rect 16865 6817 16899 6851
rect 17233 6817 17267 6851
rect 18613 6817 18647 6851
rect 1501 6749 1535 6783
rect 1961 6749 1995 6783
rect 2329 6749 2363 6783
rect 3985 6749 4019 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 7757 6749 7791 6783
rect 11161 6749 11195 6783
rect 13712 6749 13746 6783
rect 13829 6749 13863 6783
rect 13921 6749 13955 6783
rect 14381 6749 14415 6783
rect 17509 6749 17543 6783
rect 18521 6749 18555 6783
rect 3433 6681 3467 6715
rect 10057 6681 10091 6715
rect 11437 6681 11471 6715
rect 12173 6681 12207 6715
rect 13553 6681 13587 6715
rect 15669 6681 15703 6715
rect 16405 6681 16439 6715
rect 3065 6613 3099 6647
rect 3617 6613 3651 6647
rect 9413 6613 9447 6647
rect 11805 6613 11839 6647
rect 13185 6613 13219 6647
rect 4261 6409 4295 6443
rect 4997 6409 5031 6443
rect 6101 6409 6135 6443
rect 6469 6409 6503 6443
rect 11621 6409 11655 6443
rect 13645 6409 13679 6443
rect 14197 6409 14231 6443
rect 17693 6409 17727 6443
rect 18245 6409 18279 6443
rect 4859 6341 4893 6375
rect 6837 6341 6871 6375
rect 8769 6341 8803 6375
rect 11529 6341 11563 6375
rect 12633 6341 12667 6375
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 5641 6273 5675 6307
rect 7481 6273 7515 6307
rect 9229 6273 9263 6307
rect 9321 6273 9355 6307
rect 9781 6273 9815 6307
rect 10057 6273 10091 6307
rect 13277 6273 13311 6307
rect 14289 6273 14323 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 16957 6273 16991 6307
rect 18705 6273 18739 6307
rect 4537 6205 4571 6239
rect 4997 6199 5031 6233
rect 5457 6205 5491 6239
rect 5549 6205 5583 6239
rect 6193 6205 6227 6239
rect 6653 6205 6687 6239
rect 7297 6205 7331 6239
rect 8585 6205 8619 6239
rect 11805 6205 11839 6239
rect 11989 6205 12023 6239
rect 13001 6205 13035 6239
rect 13093 6205 13127 6239
rect 13369 6205 13403 6239
rect 13553 6205 13587 6239
rect 14072 6205 14106 6239
rect 15853 6205 15887 6239
rect 17049 6205 17083 6239
rect 17785 6205 17819 6239
rect 17969 6205 18003 6239
rect 18245 6205 18279 6239
rect 18429 6205 18463 6239
rect 18889 6205 18923 6239
rect 4077 6137 4111 6171
rect 4277 6137 4311 6171
rect 7205 6137 7239 6171
rect 9137 6137 9171 6171
rect 12265 6137 12299 6171
rect 12449 6137 12483 6171
rect 12817 6137 12851 6171
rect 13948 6137 13982 6171
rect 17601 6137 17635 6171
rect 4445 6069 4479 6103
rect 4629 6069 4663 6103
rect 4721 6069 4755 6103
rect 8401 6069 8435 6103
rect 19073 6069 19107 6103
rect 3985 5865 4019 5899
rect 6745 5865 6779 5899
rect 9413 5865 9447 5899
rect 10425 5865 10459 5899
rect 12633 5865 12667 5899
rect 15669 5865 15703 5899
rect 18981 5865 19015 5899
rect 2513 5797 2547 5831
rect 10977 5797 11011 5831
rect 11161 5797 11195 5831
rect 18613 5797 18647 5831
rect 2237 5729 2271 5763
rect 4353 5729 4387 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 5365 5729 5399 5763
rect 6653 5729 6687 5763
rect 7297 5729 7331 5763
rect 7665 5729 7699 5763
rect 9689 5729 9723 5763
rect 10333 5729 10367 5763
rect 11345 5729 11379 5763
rect 11529 5729 11563 5763
rect 11621 5729 11655 5763
rect 12357 5729 12391 5763
rect 12449 5729 12483 5763
rect 13461 5729 13495 5763
rect 13553 5729 13587 5763
rect 13829 5729 13863 5763
rect 14381 5729 14415 5763
rect 15761 5729 15795 5763
rect 15853 5729 15887 5763
rect 17233 5729 17267 5763
rect 17969 5729 18003 5763
rect 18889 5729 18923 5763
rect 19073 5729 19107 5763
rect 5089 5661 5123 5695
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 5825 5661 5859 5695
rect 6469 5661 6503 5695
rect 7941 5661 7975 5695
rect 10517 5661 10551 5695
rect 12081 5661 12115 5695
rect 12817 5661 12851 5695
rect 13737 5661 13771 5695
rect 14473 5661 14507 5695
rect 15485 5661 15519 5695
rect 16129 5661 16163 5695
rect 7205 5593 7239 5627
rect 9597 5593 9631 5627
rect 9965 5593 9999 5627
rect 13277 5593 13311 5627
rect 17417 5593 17451 5627
rect 4169 5525 4203 5559
rect 4905 5525 4939 5559
rect 11805 5525 11839 5559
rect 13001 5525 13035 5559
rect 3696 5321 3730 5355
rect 5457 5321 5491 5355
rect 8033 5321 8067 5355
rect 10517 5321 10551 5355
rect 16129 5321 16163 5355
rect 16865 5321 16899 5355
rect 6837 5253 6871 5287
rect 11713 5253 11747 5287
rect 15761 5253 15795 5287
rect 3433 5185 3467 5219
rect 5181 5185 5215 5219
rect 7481 5185 7515 5219
rect 8769 5185 8803 5219
rect 10977 5185 11011 5219
rect 11897 5185 11931 5219
rect 16405 5185 16439 5219
rect 18429 5185 18463 5219
rect 5733 5117 5767 5151
rect 6653 5117 6687 5151
rect 7205 5117 7239 5151
rect 10885 5117 10919 5151
rect 11161 5117 11195 5151
rect 11621 5117 11655 5151
rect 11713 5117 11747 5151
rect 12265 5117 12299 5151
rect 13369 5117 13403 5151
rect 14289 5117 14323 5151
rect 15393 5117 15427 5151
rect 15945 5117 15979 5151
rect 16313 5117 16347 5151
rect 16589 5117 16623 5151
rect 16681 5117 16715 5151
rect 16957 5117 16991 5151
rect 18521 5117 18555 5151
rect 18797 5117 18831 5151
rect 18981 5117 19015 5151
rect 7297 5049 7331 5083
rect 8125 5049 8159 5083
rect 9045 5049 9079 5083
rect 11437 5049 11471 5083
rect 13921 5049 13955 5083
rect 18705 5049 18739 5083
rect 6469 4981 6503 5015
rect 11345 4981 11379 5015
rect 13645 4981 13679 5015
rect 7757 4777 7791 4811
rect 8953 4777 8987 4811
rect 10793 4777 10827 4811
rect 11713 4777 11747 4811
rect 16221 4777 16255 4811
rect 17417 4777 17451 4811
rect 4169 4709 4203 4743
rect 6285 4709 6319 4743
rect 11069 4709 11103 4743
rect 12081 4709 12115 4743
rect 857 4641 891 4675
rect 3893 4641 3927 4675
rect 6009 4641 6043 4675
rect 8217 4641 8251 4675
rect 8309 4641 8343 4675
rect 9680 4641 9714 4675
rect 11345 4641 11379 4675
rect 14749 4641 14783 4675
rect 15853 4641 15887 4675
rect 16129 4641 16163 4675
rect 16405 4641 16439 4675
rect 16865 4641 16899 4675
rect 17141 4641 17175 4675
rect 17233 4641 17267 4675
rect 17509 4641 17543 4675
rect 19073 4641 19107 4675
rect 5641 4573 5675 4607
rect 8769 4573 8803 4607
rect 8861 4573 8895 4607
rect 9413 4573 9447 4607
rect 11253 4573 11287 4607
rect 11805 4573 11839 4607
rect 13829 4573 13863 4607
rect 16957 4573 16991 4607
rect 18521 4573 18555 4607
rect 14565 4505 14599 4539
rect 1041 4437 1075 4471
rect 8493 4437 8527 4471
rect 9321 4437 9355 4471
rect 16589 4437 16623 4471
rect 18245 4233 18279 4267
rect 9321 4165 9355 4199
rect 15393 4165 15427 4199
rect 17049 4165 17083 4199
rect 6285 4097 6319 4131
rect 8033 4097 8067 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9965 4097 9999 4131
rect 11621 4097 11655 4131
rect 11989 4097 12023 4131
rect 13369 4097 13403 4131
rect 15577 4097 15611 4131
rect 1133 4029 1167 4063
rect 1225 4029 1259 4063
rect 1409 4029 1443 4063
rect 2881 4029 2915 4063
rect 2973 4029 3007 4063
rect 3249 4029 3283 4063
rect 8769 4029 8803 4063
rect 9597 4029 9631 4063
rect 9873 4029 9907 4063
rect 10057 4029 10091 4063
rect 10149 4029 10183 4063
rect 11713 4029 11747 4063
rect 11805 4029 11839 4063
rect 13737 4029 13771 4063
rect 13921 4029 13955 4063
rect 15485 4029 15519 4063
rect 16681 4029 16715 4063
rect 18429 4029 18463 4063
rect 18889 4029 18923 4063
rect 1654 3961 1688 3995
rect 3516 3961 3550 3995
rect 6561 3961 6595 3995
rect 13645 3961 13679 3995
rect 17325 3961 17359 3995
rect 18153 3961 18187 3995
rect 2789 3893 2823 3927
rect 4629 3893 4663 3927
rect 8401 3893 8435 3927
rect 18797 3893 18831 3927
rect 3801 3689 3835 3723
rect 6745 3689 6779 3723
rect 15853 3689 15887 3723
rect 17509 3689 17543 3723
rect 11253 3621 11287 3655
rect 15117 3621 15151 3655
rect 3157 3553 3191 3587
rect 6929 3553 6963 3587
rect 9873 3553 9907 3587
rect 10149 3553 10183 3587
rect 10333 3553 10367 3587
rect 10977 3553 11011 3587
rect 13093 3553 13127 3587
rect 15209 3553 15243 3587
rect 17417 3553 17451 3587
rect 17601 3553 17635 3587
rect 18521 3553 18555 3587
rect 8125 3485 8159 3519
rect 9597 3485 9631 3519
rect 13001 3485 13035 3519
rect 13369 3485 13403 3519
rect 17969 3485 18003 3519
rect 18245 3485 18279 3519
rect 9965 3417 9999 3451
rect 10793 3417 10827 3451
rect 10609 3349 10643 3383
rect 8493 3009 8527 3043
rect 9965 3009 9999 3043
rect 10149 3009 10183 3043
rect 11437 3009 11471 3043
rect 11805 3009 11839 3043
rect 13277 3009 13311 3043
rect 13921 3009 13955 3043
rect 15117 3009 15151 3043
rect 15761 3009 15795 3043
rect 16865 3009 16899 3043
rect 18061 3009 18095 3043
rect 6837 2941 6871 2975
rect 7021 2941 7055 2975
rect 7297 2941 7331 2975
rect 7573 2941 7607 2975
rect 8217 2941 8251 2975
rect 10057 2941 10091 2975
rect 11621 2941 11655 2975
rect 12909 2941 12943 2975
rect 14013 2941 14047 2975
rect 15669 2941 15703 2975
rect 16773 2941 16807 2975
rect 17969 2941 18003 2975
rect 19073 2941 19107 2975
rect 8125 2805 8159 2839
rect 18889 2805 18923 2839
rect 18889 2601 18923 2635
rect 8002 2533 8036 2567
rect 5825 2465 5859 2499
rect 6009 2465 6043 2499
rect 6101 2465 6135 2499
rect 6285 2465 6319 2499
rect 6653 2465 6687 2499
rect 7205 2465 7239 2499
rect 7757 2465 7791 2499
rect 9229 2465 9263 2499
rect 10793 2465 10827 2499
rect 11437 2465 11471 2499
rect 12633 2465 12667 2499
rect 14105 2465 14139 2499
rect 14381 2465 14415 2499
rect 17233 2465 17267 2499
rect 18337 2465 18371 2499
rect 19073 2465 19107 2499
rect 7481 2397 7515 2431
rect 10609 2397 10643 2431
rect 11529 2397 11563 2431
rect 12541 2397 12575 2431
rect 14013 2397 14047 2431
rect 14565 2397 14599 2431
rect 15945 2397 15979 2431
rect 16129 2397 16163 2431
rect 18521 2397 18555 2431
rect 17601 2329 17635 2363
rect 6561 2261 6595 2295
rect 6929 2261 6963 2295
rect 9137 2261 9171 2295
rect 6515 2057 6549 2091
rect 8125 2057 8159 2091
rect 14013 1989 14047 2023
rect 16221 1989 16255 2023
rect 6975 1921 7009 1955
rect 8861 1921 8895 1955
rect 11621 1921 11655 1955
rect 13277 1921 13311 1955
rect 13645 1921 13679 1955
rect 16865 1921 16899 1955
rect 18061 1921 18095 1955
rect 857 1853 891 1887
rect 5733 1853 5767 1887
rect 5825 1853 5859 1887
rect 6101 1853 6135 1887
rect 6285 1853 6319 1887
rect 6444 1853 6478 1887
rect 6837 1853 6871 1887
rect 7078 1853 7112 1887
rect 7389 1853 7423 1887
rect 7481 1853 7515 1887
rect 7941 1853 7975 1887
rect 8033 1853 8067 1887
rect 8953 1853 8987 1887
rect 10057 1853 10091 1887
rect 10149 1853 10183 1887
rect 11713 1853 11747 1887
rect 11805 1853 11839 1887
rect 13369 1853 13403 1887
rect 14749 1853 14783 1887
rect 15853 1853 15887 1887
rect 17969 1853 18003 1887
rect 18889 1853 18923 1887
rect 14013 1717 14047 1751
rect 10977 1513 11011 1547
rect 15761 1445 15795 1479
rect 18521 1445 18555 1479
rect 5457 1377 5491 1411
rect 5641 1377 5675 1411
rect 6193 1377 6227 1411
rect 6377 1377 6411 1411
rect 6469 1377 6503 1411
rect 6653 1377 6687 1411
rect 6745 1377 6779 1411
rect 6929 1377 6963 1411
rect 7021 1377 7055 1411
rect 7205 1377 7239 1411
rect 7297 1377 7331 1411
rect 7481 1377 7515 1411
rect 8677 1377 8711 1411
rect 10793 1377 10827 1411
rect 11529 1377 11563 1411
rect 11713 1377 11747 1411
rect 11897 1377 11931 1411
rect 13645 1377 13679 1411
rect 14841 1377 14875 1411
rect 15485 1377 15519 1411
rect 17509 1377 17543 1411
rect 18245 1377 18279 1411
rect 19073 1377 19107 1411
rect 7573 1309 7607 1343
rect 9229 1309 9263 1343
rect 10701 1309 10735 1343
rect 12081 1309 12115 1343
rect 13737 1309 13771 1343
rect 14749 1309 14783 1343
rect 16405 1309 16439 1343
rect 17877 1309 17911 1343
rect 9045 1241 9079 1275
rect 13553 1241 13587 1275
rect 6101 1173 6135 1207
rect 8401 969 8435 1003
rect 19073 969 19107 1003
rect 8677 901 8711 935
rect 11897 901 11931 935
rect 13645 901 13679 935
rect 17601 901 17635 935
rect 6653 833 6687 867
rect 8125 833 8159 867
rect 9321 833 9355 867
rect 10793 833 10827 867
rect 13369 833 13403 867
rect 15117 833 15151 867
rect 16129 833 16163 867
rect 3985 765 4019 799
rect 5825 765 5859 799
rect 6009 765 6043 799
rect 6101 765 6135 799
rect 6285 765 6319 799
rect 6377 765 6411 799
rect 6561 765 6595 799
rect 7757 765 7791 799
rect 8953 765 8987 799
rect 9137 765 9171 799
rect 9229 765 9263 799
rect 10977 765 11011 799
rect 11161 765 11195 799
rect 11805 765 11839 799
rect 14013 765 14047 799
rect 17509 765 17543 799
rect 17785 629 17819 663
rect 18337 629 18371 663
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 3878 18912 3884 18964
rect 3936 18952 3942 18964
rect 3973 18955 4031 18961
rect 3973 18952 3985 18955
rect 3936 18924 3985 18952
rect 3936 18912 3942 18924
rect 3973 18921 3985 18924
rect 4019 18921 4031 18955
rect 3973 18915 4031 18921
rect 7742 18844 7748 18896
rect 7800 18884 7806 18896
rect 8481 18887 8539 18893
rect 8481 18884 8493 18887
rect 7800 18856 8493 18884
rect 7800 18844 7806 18856
rect 8481 18853 8493 18856
rect 8527 18853 8539 18887
rect 8481 18847 8539 18853
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 8168 18788 9413 18816
rect 8168 18776 8174 18788
rect 9401 18785 9413 18788
rect 9447 18785 9459 18819
rect 9401 18779 9459 18785
rect 15470 18776 15476 18828
rect 15528 18816 15534 18828
rect 15565 18819 15623 18825
rect 15565 18816 15577 18819
rect 15528 18788 15577 18816
rect 15528 18776 15534 18788
rect 15565 18785 15577 18788
rect 15611 18785 15623 18819
rect 15565 18779 15623 18785
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 16209 18819 16267 18825
rect 16209 18816 16221 18819
rect 16172 18788 16221 18816
rect 16172 18776 16178 18788
rect 16209 18785 16221 18788
rect 16255 18785 16267 18819
rect 16209 18779 16267 18785
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18104 18788 18153 18816
rect 18104 18776 18110 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 842 18708 848 18760
rect 900 18708 906 18760
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 9306 18708 9312 18760
rect 9364 18708 9370 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10410 18748 10416 18760
rect 9732 18720 10416 18748
rect 9732 18708 9738 18720
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 8662 18640 8668 18692
rect 8720 18640 8726 18692
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 9769 18615 9827 18621
rect 9769 18612 9781 18615
rect 9732 18584 9781 18612
rect 9732 18572 9738 18584
rect 9769 18581 9781 18584
rect 9815 18581 9827 18615
rect 9769 18575 9827 18581
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 10502 18232 10508 18284
rect 10560 18272 10566 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10560 18244 10793 18272
rect 10560 18232 10566 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 6362 18164 6368 18216
rect 6420 18164 6426 18216
rect 6086 18096 6092 18148
rect 6144 18136 6150 18148
rect 6641 18139 6699 18145
rect 6641 18136 6653 18139
rect 6144 18108 6653 18136
rect 6144 18096 6150 18108
rect 6641 18105 6653 18108
rect 6687 18105 6699 18139
rect 8938 18136 8944 18148
rect 7866 18108 8944 18136
rect 6641 18099 6699 18105
rect 8938 18096 8944 18108
rect 8996 18136 9002 18148
rect 8996 18108 9338 18136
rect 8996 18096 9002 18108
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 10505 18139 10563 18145
rect 10505 18136 10517 18139
rect 10284 18108 10517 18136
rect 10284 18096 10290 18108
rect 10505 18105 10517 18108
rect 10551 18105 10563 18139
rect 10505 18099 10563 18105
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 8110 18068 8116 18080
rect 6880 18040 8116 18068
rect 6880 18028 6886 18040
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9214 18068 9220 18080
rect 9079 18040 9220 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 7282 17864 7288 17876
rect 6840 17836 7288 17864
rect 4890 17756 4896 17808
rect 4948 17756 4954 17808
rect 6701 17799 6759 17805
rect 6701 17796 6713 17799
rect 5460 17768 6713 17796
rect 5460 17740 5488 17768
rect 6701 17765 6713 17768
rect 6747 17796 6759 17799
rect 6840 17796 6868 17836
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 9674 17824 9680 17876
rect 9732 17824 9738 17876
rect 10045 17867 10103 17873
rect 10045 17833 10057 17867
rect 10091 17864 10103 17867
rect 10226 17864 10232 17876
rect 10091 17836 10232 17864
rect 10091 17833 10103 17836
rect 10045 17827 10103 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 11149 17867 11207 17873
rect 11149 17833 11161 17867
rect 11195 17833 11207 17867
rect 11149 17827 11207 17833
rect 6747 17768 6868 17796
rect 6917 17799 6975 17805
rect 6747 17765 6759 17768
rect 6701 17759 6759 17765
rect 6917 17765 6929 17799
rect 6963 17796 6975 17799
rect 7098 17796 7104 17808
rect 6963 17768 7104 17796
rect 6963 17765 6975 17768
rect 6917 17759 6975 17765
rect 5442 17688 5448 17740
rect 5500 17688 5506 17740
rect 5629 17731 5687 17737
rect 5629 17697 5641 17731
rect 5675 17728 5687 17731
rect 5718 17728 5724 17740
rect 5675 17700 5724 17728
rect 5675 17697 5687 17700
rect 5629 17691 5687 17697
rect 5718 17688 5724 17700
rect 5776 17728 5782 17740
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 5776 17700 6469 17728
rect 5776 17688 5782 17700
rect 6457 17697 6469 17700
rect 6503 17728 6515 17731
rect 6932 17728 6960 17759
rect 7098 17756 7104 17768
rect 7156 17756 7162 17808
rect 7374 17756 7380 17808
rect 7432 17796 7438 17808
rect 7469 17799 7527 17805
rect 7469 17796 7481 17799
rect 7432 17768 7481 17796
rect 7432 17756 7438 17768
rect 7469 17765 7481 17768
rect 7515 17765 7527 17799
rect 7469 17759 7527 17765
rect 8938 17728 8944 17740
rect 6503 17700 6960 17728
rect 8602 17700 8944 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9692 17728 9720 17824
rect 11164 17796 11192 17827
rect 11517 17799 11575 17805
rect 11517 17796 11529 17799
rect 11164 17768 11529 17796
rect 11517 17765 11529 17768
rect 11563 17765 11575 17799
rect 11517 17759 11575 17765
rect 12526 17756 12532 17808
rect 12584 17756 12590 17808
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9692 17700 9873 17728
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10962 17688 10968 17740
rect 11020 17688 11026 17740
rect 3510 17620 3516 17672
rect 3568 17660 3574 17672
rect 3605 17663 3663 17669
rect 3605 17660 3617 17663
rect 3568 17632 3617 17660
rect 3568 17620 3574 17632
rect 3605 17629 3617 17632
rect 3651 17629 3663 17663
rect 3605 17623 3663 17629
rect 3878 17620 3884 17672
rect 3936 17620 3942 17672
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 6420 17632 7205 17660
rect 6420 17620 6426 17632
rect 7193 17629 7205 17632
rect 7239 17660 7251 17663
rect 8846 17660 8852 17672
rect 7239 17632 8852 17660
rect 7239 17629 7251 17632
rect 7193 17623 7251 17629
rect 8846 17620 8852 17632
rect 8904 17620 8910 17672
rect 10502 17620 10508 17672
rect 10560 17660 10566 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 10560 17632 11253 17660
rect 10560 17620 10566 17632
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 5810 17484 5816 17536
rect 5868 17484 5874 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 6549 17527 6607 17533
rect 6549 17524 6561 17527
rect 6420 17496 6561 17524
rect 6420 17484 6426 17496
rect 6549 17493 6561 17496
rect 6595 17493 6607 17527
rect 6549 17487 6607 17493
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 6822 17524 6828 17536
rect 6779 17496 6828 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 8941 17527 8999 17533
rect 8941 17524 8953 17527
rect 7248 17496 8953 17524
rect 7248 17484 7254 17496
rect 8941 17493 8953 17496
rect 8987 17524 8999 17527
rect 11882 17524 11888 17536
rect 8987 17496 11888 17524
rect 8987 17493 8999 17496
rect 8941 17487 8999 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12676 17496 13001 17524
rect 12676 17484 12682 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 3878 17280 3884 17332
rect 3936 17320 3942 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 3936 17292 4445 17320
rect 3936 17280 3942 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 4801 17323 4859 17329
rect 4801 17289 4813 17323
rect 4847 17320 4859 17323
rect 4847 17292 5488 17320
rect 4847 17289 4859 17292
rect 4801 17283 4859 17289
rect 5460 17264 5488 17292
rect 5810 17280 5816 17332
rect 5868 17280 5874 17332
rect 6086 17280 6092 17332
rect 6144 17280 6150 17332
rect 7285 17323 7343 17329
rect 6288 17292 7236 17320
rect 4985 17255 5043 17261
rect 4985 17221 4997 17255
rect 5031 17221 5043 17255
rect 4985 17215 5043 17221
rect 5000 17184 5028 17215
rect 5442 17212 5448 17264
rect 5500 17212 5506 17264
rect 5828 17184 5856 17280
rect 6181 17255 6239 17261
rect 6181 17221 6193 17255
rect 6227 17252 6239 17255
rect 6288 17252 6316 17292
rect 6227 17224 6316 17252
rect 6227 17221 6239 17224
rect 6181 17215 6239 17221
rect 6362 17212 6368 17264
rect 6420 17252 6426 17264
rect 7208 17252 7236 17292
rect 7285 17289 7297 17323
rect 7331 17320 7343 17323
rect 7374 17320 7380 17332
rect 7331 17292 7380 17320
rect 7331 17289 7343 17292
rect 7285 17283 7343 17289
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 11425 17323 11483 17329
rect 11425 17320 11437 17323
rect 11020 17292 11437 17320
rect 11020 17280 11026 17292
rect 11425 17289 11437 17292
rect 11471 17289 11483 17323
rect 11425 17283 11483 17289
rect 7653 17255 7711 17261
rect 7653 17252 7665 17255
rect 6420 17224 6960 17252
rect 7208 17224 7665 17252
rect 6420 17212 6426 17224
rect 6457 17187 6515 17193
rect 4632 17156 5028 17184
rect 5184 17156 5856 17184
rect 6104 17156 6408 17184
rect 4632 17125 4660 17156
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17116 4951 17119
rect 5184 17116 5212 17156
rect 4939 17088 5212 17116
rect 5261 17119 5319 17125
rect 4939 17085 4951 17088
rect 4893 17079 4951 17085
rect 5261 17085 5273 17119
rect 5307 17116 5319 17119
rect 5442 17116 5448 17128
rect 5307 17088 5448 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 5442 17076 5448 17088
rect 5500 17116 5506 17128
rect 6104 17116 6132 17156
rect 5500 17088 6132 17116
rect 5500 17076 5506 17088
rect 6270 17076 6276 17128
rect 6328 17076 6334 17128
rect 6380 17125 6408 17156
rect 6457 17153 6469 17187
rect 6503 17184 6515 17187
rect 6503 17156 6868 17184
rect 6503 17153 6515 17156
rect 6457 17147 6515 17153
rect 6365 17119 6423 17125
rect 6365 17085 6377 17119
rect 6411 17085 6423 17119
rect 6365 17079 6423 17085
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 4985 17051 5043 17057
rect 4985 17017 4997 17051
rect 5031 17048 5043 17051
rect 5534 17048 5540 17060
rect 5031 17020 5540 17048
rect 5031 17017 5043 17020
rect 4985 17011 5043 17017
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 5626 17008 5632 17060
rect 5684 17048 5690 17060
rect 5997 17051 6055 17057
rect 5997 17048 6009 17051
rect 5684 17020 6009 17048
rect 5684 17008 5690 17020
rect 5997 17017 6009 17020
rect 6043 17017 6055 17051
rect 6564 17048 6592 17079
rect 6638 17076 6644 17128
rect 6696 17076 6702 17128
rect 6840 17125 6868 17156
rect 6932 17125 6960 17224
rect 7653 17221 7665 17224
rect 7699 17221 7711 17255
rect 7653 17215 7711 17221
rect 7098 17144 7104 17196
rect 7156 17184 7162 17196
rect 10502 17184 10508 17196
rect 7156 17156 7512 17184
rect 7156 17144 7162 17156
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7055 17088 7236 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 6564 17020 7144 17048
rect 5997 17011 6055 17017
rect 7116 16992 7144 17020
rect 7208 16992 7236 17088
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 7340 17088 7389 17116
rect 7340 17076 7346 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 5718 16980 5724 16992
rect 5215 16952 5724 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 7098 16940 7104 16992
rect 7156 16940 7162 16992
rect 7190 16940 7196 16992
rect 7248 16940 7254 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7484 16989 7512 17156
rect 9048 17156 10508 17184
rect 8754 17076 8760 17128
rect 8812 17076 8818 17128
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 9048 17125 9076 17156
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11756 17156 11989 17184
rect 11756 17144 11762 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 9033 17119 9091 17125
rect 9033 17116 9045 17119
rect 8904 17088 9045 17116
rect 8904 17076 8910 17088
rect 9033 17085 9045 17088
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 11885 17119 11943 17125
rect 11885 17085 11897 17119
rect 11931 17116 11943 17119
rect 12618 17116 12624 17128
rect 11931 17088 12624 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 7653 17051 7711 17057
rect 7653 17048 7665 17051
rect 7616 17020 7665 17048
rect 7616 17008 7622 17020
rect 7653 17017 7665 17020
rect 7699 17017 7711 17051
rect 9309 17051 9367 17057
rect 9309 17048 9321 17051
rect 7653 17011 7711 17017
rect 8956 17020 9321 17048
rect 8956 16989 8984 17020
rect 9309 17017 9321 17020
rect 9355 17017 9367 17051
rect 12526 17048 12532 17060
rect 10534 17020 12532 17048
rect 9309 17011 9367 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 7469 16983 7527 16989
rect 7469 16980 7481 16983
rect 7432 16952 7481 16980
rect 7432 16940 7438 16952
rect 7469 16949 7481 16952
rect 7515 16949 7527 16983
rect 7469 16943 7527 16949
rect 8941 16983 8999 16989
rect 8941 16949 8953 16983
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 10594 16980 10600 16992
rect 9732 16952 10600 16980
rect 9732 16940 9738 16952
rect 10594 16940 10600 16952
rect 10652 16980 10658 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10652 16952 10793 16980
rect 10652 16940 10658 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 11793 16983 11851 16989
rect 11793 16949 11805 16983
rect 11839 16980 11851 16983
rect 11882 16980 11888 16992
rect 11839 16952 11888 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 6696 16748 7052 16776
rect 6696 16736 6702 16748
rect 6914 16708 6920 16720
rect 6656 16680 6920 16708
rect 3694 16600 3700 16652
rect 3752 16600 3758 16652
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5534 16640 5540 16652
rect 5307 16612 5540 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5534 16600 5540 16612
rect 5592 16640 5598 16652
rect 6178 16640 6184 16652
rect 5592 16612 6184 16640
rect 5592 16600 5598 16612
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6656 16649 6684 16680
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 6730 16600 6736 16652
rect 6788 16600 6794 16652
rect 7024 16649 7052 16748
rect 7098 16736 7104 16788
rect 7156 16736 7162 16788
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 8754 16776 8760 16788
rect 8619 16748 8760 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 9033 16779 9091 16785
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9674 16776 9680 16788
rect 9079 16748 9680 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 7248 16677 7312 16708
rect 7248 16668 7251 16677
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16609 7067 16643
rect 7239 16643 7251 16668
rect 7285 16646 7312 16677
rect 7374 16668 7380 16720
rect 7432 16708 7438 16720
rect 7469 16711 7527 16717
rect 7469 16708 7481 16711
rect 7432 16680 7481 16708
rect 7432 16668 7438 16680
rect 7469 16677 7481 16680
rect 7515 16708 7527 16711
rect 8941 16711 8999 16717
rect 8941 16708 8953 16711
rect 7515 16680 8953 16708
rect 7515 16677 7527 16680
rect 7469 16671 7527 16677
rect 8941 16677 8953 16680
rect 8987 16677 8999 16711
rect 8941 16671 8999 16677
rect 7285 16643 7297 16646
rect 7239 16637 7297 16643
rect 7009 16603 7067 16609
rect 5902 16532 5908 16584
rect 5960 16572 5966 16584
rect 6840 16572 6868 16603
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 18785 16643 18843 16649
rect 18785 16640 18797 16643
rect 15804 16612 18797 16640
rect 15804 16600 15810 16612
rect 18785 16609 18797 16612
rect 18831 16609 18843 16643
rect 18785 16603 18843 16609
rect 18966 16600 18972 16652
rect 19024 16600 19030 16652
rect 5960 16544 6868 16572
rect 5960 16532 5966 16544
rect 9122 16532 9128 16584
rect 9180 16532 9186 16584
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 3513 16439 3571 16445
rect 3513 16436 3525 16439
rect 3476 16408 3525 16436
rect 3476 16396 3482 16408
rect 3513 16405 3525 16408
rect 3559 16405 3571 16439
rect 3513 16399 3571 16405
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 6362 16396 6368 16448
rect 6420 16396 6426 16448
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 7285 16439 7343 16445
rect 7285 16436 7297 16439
rect 6880 16408 7297 16436
rect 6880 16396 6886 16408
rect 7285 16405 7297 16408
rect 7331 16436 7343 16439
rect 7558 16436 7564 16448
rect 7331 16408 7564 16436
rect 7331 16405 7343 16408
rect 7285 16399 7343 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 6638 16232 6644 16244
rect 4028 16204 6644 16232
rect 4028 16192 4034 16204
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 6972 16204 7297 16232
rect 6972 16192 6978 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 7285 16195 7343 16201
rect 7392 16204 11560 16232
rect 4982 16124 4988 16176
rect 5040 16164 5046 16176
rect 7392 16164 7420 16204
rect 5040 16136 7420 16164
rect 8864 16136 9674 16164
rect 5040 16124 5046 16136
rect 8864 16108 8892 16136
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16096 3295 16099
rect 3510 16096 3516 16108
rect 3283 16068 3516 16096
rect 3283 16065 3295 16068
rect 3237 16059 3295 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9122 16096 9128 16108
rect 9079 16068 9128 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9646 16096 9674 16136
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9646 16068 9873 16096
rect 9861 16065 9873 16068
rect 9907 16096 9919 16099
rect 11422 16096 11428 16108
rect 9907 16068 11428 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 7193 16031 7251 16037
rect 3418 15920 3424 15972
rect 3476 15960 3482 15972
rect 3513 15963 3571 15969
rect 3513 15960 3525 15963
rect 3476 15932 3525 15960
rect 3476 15920 3482 15932
rect 3513 15929 3525 15932
rect 3559 15929 3571 15963
rect 3513 15923 3571 15929
rect 4338 15852 4344 15904
rect 4396 15892 4402 15904
rect 4632 15892 4660 16014
rect 7193 15997 7205 16031
rect 7239 16028 7251 16031
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7239 16000 7849 16028
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 7852 15904 7880 15991
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 11532 15972 11560 16204
rect 12437 16167 12495 16173
rect 12437 16133 12449 16167
rect 12483 16133 12495 16167
rect 12437 16127 12495 16133
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 11756 16068 11805 16096
rect 11756 16056 11762 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12066 16028 12072 16040
rect 12023 16000 12072 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 12452 16028 12480 16127
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12452 16000 12725 16028
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 19058 16028 19064 16040
rect 19015 16000 19064 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 9784 15932 10149 15960
rect 4396 15864 4660 15892
rect 4396 15852 4402 15864
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 5776 15864 6561 15892
rect 5776 15852 5782 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6549 15855 6607 15861
rect 7834 15852 7840 15904
rect 7892 15852 7898 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 8352 15864 8401 15892
rect 8352 15852 8358 15864
rect 8389 15861 8401 15864
rect 8435 15861 8447 15895
rect 8389 15855 8447 15861
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 8757 15895 8815 15901
rect 8757 15892 8769 15895
rect 8536 15864 8769 15892
rect 8536 15852 8542 15864
rect 8757 15861 8769 15864
rect 8803 15861 8815 15895
rect 8757 15855 8815 15861
rect 8849 15895 8907 15901
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 9214 15892 9220 15904
rect 8895 15864 9220 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 9784 15901 9812 15932
rect 10137 15929 10149 15932
rect 10183 15929 10195 15963
rect 10137 15923 10195 15929
rect 10686 15920 10692 15972
rect 10744 15920 10750 15972
rect 11514 15920 11520 15972
rect 11572 15960 11578 15972
rect 11572 15932 12112 15960
rect 11572 15920 11578 15932
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15861 9827 15895
rect 9769 15855 9827 15861
rect 11606 15852 11612 15904
rect 11664 15852 11670 15904
rect 12084 15901 12112 15932
rect 12069 15895 12127 15901
rect 12069 15861 12081 15895
rect 12115 15861 12127 15895
rect 12069 15855 12127 15861
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12308 15864 12541 15892
rect 12308 15852 12314 15864
rect 12529 15861 12541 15864
rect 12575 15861 12587 15895
rect 12529 15855 12587 15861
rect 16574 15852 16580 15904
rect 16632 15892 16638 15904
rect 18785 15895 18843 15901
rect 18785 15892 18797 15895
rect 16632 15864 18797 15892
rect 16632 15852 16638 15864
rect 18785 15861 18797 15864
rect 18831 15861 18843 15895
rect 18785 15855 18843 15861
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 5442 15688 5448 15700
rect 4632 15660 5448 15688
rect 3773 15623 3831 15629
rect 3773 15589 3785 15623
rect 3819 15620 3831 15623
rect 3878 15620 3884 15632
rect 3819 15592 3884 15620
rect 3819 15589 3831 15592
rect 3773 15583 3831 15589
rect 3878 15580 3884 15592
rect 3936 15580 3942 15632
rect 3970 15580 3976 15632
rect 4028 15580 4034 15632
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15552 2927 15555
rect 3142 15552 3148 15564
rect 2915 15524 3148 15552
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 3142 15512 3148 15524
rect 3200 15552 3206 15564
rect 4341 15555 4399 15561
rect 3200 15524 4108 15552
rect 3200 15512 3206 15524
rect 3694 15444 3700 15496
rect 3752 15444 3758 15496
rect 3605 15419 3663 15425
rect 3605 15385 3617 15419
rect 3651 15416 3663 15419
rect 3712 15416 3740 15444
rect 4080 15428 4108 15524
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4632 15552 4660 15660
rect 5442 15648 5448 15660
rect 5500 15688 5506 15700
rect 5500 15660 5856 15688
rect 5500 15648 5506 15660
rect 5718 15620 5724 15632
rect 5460 15592 5724 15620
rect 5460 15561 5488 15592
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 4387 15524 4660 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4632 15496 4660 15524
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 5626 15552 5632 15564
rect 5583 15524 5632 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 5828 15561 5856 15660
rect 5902 15648 5908 15700
rect 5960 15648 5966 15700
rect 6104 15660 7972 15688
rect 6104 15564 6132 15660
rect 6362 15580 6368 15632
rect 6420 15580 6426 15632
rect 7944 15564 7972 15660
rect 9122 15648 9128 15700
rect 9180 15688 9186 15700
rect 9180 15660 9536 15688
rect 9180 15648 9186 15660
rect 8202 15580 8208 15632
rect 8260 15580 8266 15632
rect 8938 15580 8944 15632
rect 8996 15580 9002 15632
rect 9508 15620 9536 15660
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9640 15660 9965 15688
rect 9640 15648 9646 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 9953 15651 10011 15657
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 11238 15688 11244 15700
rect 10459 15660 11244 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 11238 15648 11244 15660
rect 11296 15688 11302 15700
rect 11606 15688 11612 15700
rect 11296 15660 11612 15688
rect 11296 15648 11302 15660
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 11698 15648 11704 15700
rect 11756 15648 11762 15700
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12124 15660 13461 15688
rect 12124 15648 12130 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 11716 15620 11744 15648
rect 9508 15592 11744 15620
rect 11977 15623 12035 15629
rect 9646 15564 9674 15592
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 5994 15512 6000 15564
rect 6052 15512 6058 15564
rect 6086 15512 6092 15564
rect 6144 15512 6150 15564
rect 4614 15444 4620 15496
rect 4672 15444 4678 15496
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5353 15487 5411 15493
rect 5353 15453 5365 15487
rect 5399 15484 5411 15487
rect 5902 15484 5908 15496
rect 5399 15456 5908 15484
rect 5399 15453 5411 15456
rect 5353 15447 5411 15453
rect 3651 15388 3740 15416
rect 3651 15385 3663 15388
rect 3605 15379 3663 15385
rect 4062 15376 4068 15428
rect 4120 15376 4126 15428
rect 5276 15416 5304 15447
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 6730 15484 6736 15496
rect 6012 15456 6736 15484
rect 6012 15416 6040 15456
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 7484 15484 7512 15538
rect 7926 15512 7932 15564
rect 7984 15512 7990 15564
rect 9582 15512 9588 15564
rect 9640 15524 9674 15564
rect 9640 15512 9646 15524
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10284 15524 10333 15552
rect 10284 15512 10290 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 8938 15484 8944 15496
rect 7484 15456 8944 15484
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9677 15487 9735 15493
rect 9677 15484 9689 15487
rect 9272 15456 9689 15484
rect 9272 15444 9278 15456
rect 9677 15453 9689 15456
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 5276 15388 6040 15416
rect 1854 15308 1860 15360
rect 1912 15348 1918 15360
rect 2317 15351 2375 15357
rect 2317 15348 2329 15351
rect 1912 15320 2329 15348
rect 1912 15308 1918 15320
rect 2317 15317 2329 15320
rect 2363 15317 2375 15351
rect 2317 15311 2375 15317
rect 3789 15351 3847 15357
rect 3789 15317 3801 15351
rect 3835 15348 3847 15351
rect 4249 15351 4307 15357
rect 4249 15348 4261 15351
rect 3835 15320 4261 15348
rect 3835 15317 3847 15320
rect 3789 15311 3847 15317
rect 4249 15317 4261 15320
rect 4295 15317 4307 15351
rect 4249 15311 4307 15317
rect 5077 15351 5135 15357
rect 5077 15317 5089 15351
rect 5123 15348 5135 15351
rect 5166 15348 5172 15360
rect 5123 15320 5172 15348
rect 5123 15317 5135 15320
rect 5077 15311 5135 15317
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 6546 15308 6552 15360
rect 6604 15348 6610 15360
rect 7834 15348 7840 15360
rect 6604 15320 7840 15348
rect 6604 15308 6610 15320
rect 7834 15308 7840 15320
rect 7892 15348 7898 15360
rect 10244 15348 10272 15512
rect 10520 15493 10548 15592
rect 11977 15589 11989 15623
rect 12023 15620 12035 15623
rect 12250 15620 12256 15632
rect 12023 15592 12256 15620
rect 12023 15589 12035 15592
rect 11977 15583 12035 15589
rect 12250 15580 12256 15592
rect 12308 15580 12314 15632
rect 12526 15580 12532 15632
rect 12584 15580 12590 15632
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 11480 15524 11713 15552
rect 11480 15512 11486 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 17494 15444 17500 15496
rect 17552 15444 17558 15496
rect 18322 15444 18328 15496
rect 18380 15484 18386 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18380 15456 18521 15484
rect 18380 15444 18386 15456
rect 18509 15453 18521 15456
rect 18555 15484 18567 15487
rect 18616 15484 18644 15515
rect 18555 15456 18644 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 7892 15320 10272 15348
rect 7892 15308 7898 15320
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 3878 15104 3884 15156
rect 3936 15104 3942 15156
rect 4614 15104 4620 15156
rect 4672 15104 4678 15156
rect 4890 15104 4896 15156
rect 4948 15144 4954 15156
rect 4948 15116 6316 15144
rect 4948 15104 4954 15116
rect 3528 15076 3556 15104
rect 4798 15076 4804 15088
rect 3528 15048 4804 15076
rect 4798 15036 4804 15048
rect 4856 15076 4862 15088
rect 4856 15048 5028 15076
rect 4856 15036 4862 15048
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3142 15008 3148 15020
rect 2924 14980 3148 15008
rect 2924 14968 2930 14980
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 15008 3571 15011
rect 3970 15008 3976 15020
rect 3559 14980 3976 15008
rect 3559 14977 3571 14980
rect 3513 14971 3571 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 5000 15017 5028 15048
rect 4985 15011 5043 15017
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 842 14900 848 14952
rect 900 14900 906 14952
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3329 14943 3387 14949
rect 3329 14909 3341 14943
rect 3375 14940 3387 14943
rect 3418 14940 3424 14952
rect 3375 14912 3424 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 1118 14832 1124 14884
rect 1176 14832 1182 14884
rect 2682 14872 2688 14884
rect 2346 14844 2688 14872
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 3252 14872 3280 14903
rect 3418 14900 3424 14912
rect 3476 14940 3482 14952
rect 4062 14940 4068 14952
rect 3476 14912 4068 14940
rect 3476 14900 3482 14912
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4154 14900 4160 14952
rect 4212 14900 4218 14952
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 4890 14940 4896 14952
rect 4847 14912 4896 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 4264 14872 4292 14900
rect 3252 14844 4292 14872
rect 4356 14872 4384 14903
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 6288 14940 6316 15116
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 6788 15116 6837 15144
rect 6788 15104 6794 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 7006 15104 7012 15156
rect 7064 15104 7070 15156
rect 8202 15104 8208 15156
rect 8260 15104 8266 15156
rect 8478 15076 8484 15088
rect 6748 15048 8484 15076
rect 6748 15020 6776 15048
rect 8478 15036 8484 15048
rect 8536 15036 8542 15088
rect 8757 15079 8815 15085
rect 8757 15045 8769 15079
rect 8803 15076 8815 15079
rect 8938 15076 8944 15088
rect 8803 15048 8944 15076
rect 8803 15045 8815 15048
rect 8757 15039 8815 15045
rect 8938 15036 8944 15048
rect 8996 15076 9002 15088
rect 8996 15048 9260 15076
rect 8996 15036 9002 15048
rect 6730 14968 6736 15020
rect 6788 14968 6794 15020
rect 9232 15008 9260 15048
rect 18322 15036 18328 15088
rect 18380 15036 18386 15088
rect 12526 15008 12532 15020
rect 6840 14980 7328 15008
rect 9232 14980 12532 15008
rect 6840 14940 6868 14980
rect 6288 14912 6868 14940
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 6972 14912 7236 14940
rect 6972 14900 6978 14912
rect 4982 14872 4988 14884
rect 4356 14844 4988 14872
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 5166 14832 5172 14884
rect 5224 14872 5230 14884
rect 7208 14881 7236 14912
rect 7300 14884 7328 14980
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8294 14940 8300 14952
rect 8067 14912 8300 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8938 14900 8944 14952
rect 8996 14940 9002 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8996 14912 9137 14940
rect 8996 14900 9002 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 10520 14926 10548 14980
rect 12526 14968 12532 14980
rect 12584 15008 12590 15020
rect 16853 15011 16911 15017
rect 12584 14980 13032 15008
rect 12584 14968 12590 14980
rect 9125 14903 9183 14909
rect 11330 14900 11336 14952
rect 11388 14900 11394 14952
rect 11422 14900 11428 14952
rect 11480 14940 11486 14952
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11480 14912 11621 14940
rect 11480 14900 11486 14912
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 13004 14926 13032 14980
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 16942 15008 16948 15020
rect 16899 14980 16948 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 16942 14968 16948 14980
rect 17000 15008 17006 15020
rect 17494 15008 17500 15020
rect 17000 14980 17500 15008
rect 17000 14968 17006 14980
rect 17494 14968 17500 14980
rect 17552 14968 17558 15020
rect 18340 14949 18368 15036
rect 18325 14943 18383 14949
rect 11609 14903 11667 14909
rect 18325 14909 18337 14943
rect 18371 14909 18383 14943
rect 18325 14903 18383 14909
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 5224 14844 5273 14872
rect 5224 14832 5230 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14841 7251 14875
rect 7193 14835 7251 14841
rect 7282 14832 7288 14884
rect 7340 14872 7346 14884
rect 8481 14875 8539 14881
rect 8481 14872 8493 14875
rect 7340 14844 8493 14872
rect 7340 14832 7346 14844
rect 8481 14841 8493 14844
rect 8527 14841 8539 14875
rect 8481 14835 8539 14841
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3513 14807 3571 14813
rect 3513 14804 3525 14807
rect 3200 14776 3525 14804
rect 3200 14764 3206 14776
rect 3513 14773 3525 14776
rect 3559 14773 3571 14807
rect 3513 14767 3571 14773
rect 6993 14807 7051 14813
rect 6993 14773 7005 14807
rect 7039 14804 7051 14807
rect 7098 14804 7104 14816
rect 7039 14776 7104 14804
rect 7039 14773 7051 14776
rect 6993 14767 7051 14773
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 8496 14804 8524 14835
rect 9398 14832 9404 14884
rect 9456 14832 9462 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11532 14844 11897 14872
rect 10686 14804 10692 14816
rect 8496 14776 10692 14804
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 11532 14813 11560 14844
rect 11885 14841 11897 14844
rect 11931 14841 11943 14875
rect 11885 14835 11943 14841
rect 15838 14832 15844 14884
rect 15896 14872 15902 14884
rect 18785 14875 18843 14881
rect 18785 14872 18797 14875
rect 15896 14844 18797 14872
rect 15896 14832 15902 14844
rect 18785 14841 18797 14844
rect 18831 14841 18843 14875
rect 18785 14835 18843 14841
rect 18969 14875 19027 14881
rect 18969 14841 18981 14875
rect 19015 14872 19027 14875
rect 19058 14872 19064 14884
rect 19015 14844 19064 14872
rect 19015 14841 19027 14844
rect 18969 14835 19027 14841
rect 19058 14832 19064 14844
rect 19116 14832 19122 14884
rect 11517 14807 11575 14813
rect 11517 14773 11529 14807
rect 11563 14773 11575 14807
rect 11517 14767 11575 14773
rect 13354 14764 13360 14816
rect 13412 14764 13418 14816
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 1118 14560 1124 14612
rect 1176 14600 1182 14612
rect 1397 14603 1455 14609
rect 1397 14600 1409 14603
rect 1176 14572 1409 14600
rect 1176 14560 1182 14572
rect 1397 14569 1409 14572
rect 1443 14569 1455 14603
rect 1397 14563 1455 14569
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2179 14572 2360 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2332 14532 2360 14572
rect 2406 14560 2412 14612
rect 2464 14600 2470 14612
rect 3510 14600 3516 14612
rect 2464 14572 3516 14600
rect 2464 14560 2470 14572
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 4120 14572 4629 14600
rect 4120 14560 4126 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 4801 14603 4859 14609
rect 4801 14569 4813 14603
rect 4847 14600 4859 14603
rect 4890 14600 4896 14612
rect 4847 14572 4896 14600
rect 4847 14569 4859 14572
rect 4801 14563 4859 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 6181 14603 6239 14609
rect 6181 14600 6193 14603
rect 5500 14572 6193 14600
rect 5500 14560 5506 14572
rect 6181 14569 6193 14572
rect 6227 14600 6239 14603
rect 7006 14600 7012 14612
rect 6227 14572 7012 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8938 14600 8944 14612
rect 7984 14572 8944 14600
rect 7984 14560 7990 14572
rect 8938 14560 8944 14572
rect 8996 14600 9002 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8996 14572 9045 14600
rect 8996 14560 9002 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 9398 14560 9404 14612
rect 9456 14600 9462 14612
rect 9585 14603 9643 14609
rect 9585 14600 9597 14603
rect 9456 14572 9597 14600
rect 9456 14560 9462 14572
rect 9585 14569 9597 14572
rect 9631 14569 9643 14603
rect 9585 14563 9643 14569
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 11388 14572 11713 14600
rect 11388 14560 11394 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 11701 14563 11759 14569
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 14976 14572 16528 14600
rect 14976 14560 14982 14572
rect 2866 14532 2872 14544
rect 2332 14504 2872 14532
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4433 14535 4491 14541
rect 4433 14532 4445 14535
rect 4212 14504 4445 14532
rect 4212 14492 4218 14504
rect 4433 14501 4445 14504
rect 4479 14532 4491 14535
rect 4479 14504 5488 14532
rect 4479 14501 4491 14504
rect 4433 14495 4491 14501
rect 5460 14476 5488 14504
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 5813 14535 5871 14541
rect 5813 14532 5825 14535
rect 5684 14504 5825 14532
rect 5684 14492 5690 14504
rect 5813 14501 5825 14504
rect 5859 14501 5871 14535
rect 5813 14495 5871 14501
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 6273 14535 6331 14541
rect 6273 14532 6285 14535
rect 6052 14504 6285 14532
rect 6052 14492 6058 14504
rect 6273 14501 6285 14504
rect 6319 14501 6331 14535
rect 6273 14495 6331 14501
rect 6730 14492 6736 14544
rect 6788 14492 6794 14544
rect 15010 14492 15016 14544
rect 15068 14532 15074 14544
rect 16500 14532 16528 14572
rect 16574 14532 16580 14544
rect 15068 14504 16344 14532
rect 15068 14492 15074 14504
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1627 14436 1716 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 1688 14328 1716 14436
rect 1854 14424 1860 14476
rect 1912 14424 1918 14476
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2038 14464 2044 14476
rect 1995 14436 2044 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 2148 14436 2237 14464
rect 2148 14408 2176 14436
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 2225 14427 2283 14433
rect 2314 14424 2320 14476
rect 2372 14424 2378 14476
rect 4338 14464 4344 14476
rect 3726 14450 4344 14464
rect 3712 14436 4344 14450
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 2130 14396 2136 14408
rect 1811 14368 2136 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 1949 14331 2007 14337
rect 1949 14328 1961 14331
rect 1688 14300 1961 14328
rect 1949 14297 1961 14300
rect 1995 14297 2007 14331
rect 1949 14291 2007 14297
rect 842 14220 848 14272
rect 900 14260 906 14272
rect 2332 14260 2360 14424
rect 2590 14356 2596 14408
rect 2648 14356 2654 14408
rect 2682 14356 2688 14408
rect 2740 14396 2746 14408
rect 3712 14396 3740 14436
rect 4338 14424 4344 14436
rect 4396 14424 4402 14476
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 4982 14464 4988 14476
rect 4571 14436 4988 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 6549 14467 6607 14473
rect 5500 14436 6040 14464
rect 5500 14424 5506 14436
rect 2740 14368 3740 14396
rect 5905 14399 5963 14405
rect 2740 14356 2746 14368
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 6012 14396 6040 14436
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 6748 14464 6776 14492
rect 6595 14436 6776 14464
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7064 14436 7757 14464
rect 7064 14424 7070 14436
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 9769 14467 9827 14473
rect 9769 14464 9781 14467
rect 9732 14436 9781 14464
rect 9732 14424 9738 14436
rect 9769 14433 9781 14436
rect 9815 14433 9827 14467
rect 11974 14464 11980 14476
rect 9769 14427 9827 14433
rect 9876 14436 11980 14464
rect 9876 14396 9904 14436
rect 11974 14424 11980 14436
rect 12032 14464 12038 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 12032 14436 12081 14464
rect 12032 14424 12038 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12161 14467 12219 14473
rect 12161 14433 12173 14467
rect 12207 14464 12219 14467
rect 13078 14464 13084 14476
rect 12207 14436 13084 14464
rect 12207 14433 12219 14436
rect 12161 14427 12219 14433
rect 13078 14424 13084 14436
rect 13136 14464 13142 14476
rect 13354 14464 13360 14476
rect 13136 14436 13360 14464
rect 13136 14424 13142 14436
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 14369 14467 14427 14473
rect 14369 14433 14381 14467
rect 14415 14464 14427 14467
rect 15105 14467 15163 14473
rect 14415 14436 15056 14464
rect 14415 14433 14427 14436
rect 14369 14427 14427 14433
rect 6012 14368 9904 14396
rect 5905 14359 5963 14365
rect 4065 14331 4123 14337
rect 4065 14297 4077 14331
rect 4111 14328 4123 14331
rect 4246 14328 4252 14340
rect 4111 14300 4252 14328
rect 4111 14297 4123 14300
rect 4065 14291 4123 14297
rect 4246 14288 4252 14300
rect 4304 14288 4310 14340
rect 5920 14328 5948 14359
rect 11698 14356 11704 14408
rect 11756 14396 11762 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 11756 14368 12265 14396
rect 11756 14356 11762 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 12584 14368 14565 14396
rect 12584 14356 12590 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 15028 14396 15056 14436
rect 15105 14433 15117 14467
rect 15151 14464 15163 14467
rect 15286 14464 15292 14476
rect 15151 14436 15292 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 15286 14424 15292 14436
rect 15344 14464 15350 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15344 14436 15577 14464
rect 15344 14424 15350 14436
rect 15565 14433 15577 14436
rect 15611 14464 15623 14467
rect 15838 14464 15844 14476
rect 15611 14436 15844 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 16316 14473 16344 14504
rect 16500 14504 16580 14532
rect 16500 14473 16528 14504
rect 16574 14492 16580 14504
rect 16632 14532 16638 14544
rect 16632 14504 17356 14532
rect 16632 14492 16638 14504
rect 17328 14476 17356 14504
rect 16301 14467 16359 14473
rect 16301 14433 16313 14467
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14464 16911 14467
rect 16899 14436 17080 14464
rect 16899 14433 16911 14436
rect 16853 14427 16911 14433
rect 15194 14396 15200 14408
rect 15028 14368 15200 14396
rect 14553 14359 14611 14365
rect 15194 14356 15200 14368
rect 15252 14396 15258 14408
rect 15746 14396 15752 14408
rect 15252 14368 15752 14396
rect 15252 14356 15258 14368
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14365 16175 14399
rect 16316 14396 16344 14427
rect 16868 14396 16896 14427
rect 16316 14368 16896 14396
rect 16117 14359 16175 14365
rect 6178 14328 6184 14340
rect 5920 14300 6184 14328
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 10134 14288 10140 14340
rect 10192 14328 10198 14340
rect 10686 14328 10692 14340
rect 10192 14300 10692 14328
rect 10192 14288 10198 14300
rect 10686 14288 10692 14300
rect 10744 14328 10750 14340
rect 10870 14328 10876 14340
rect 10744 14300 10876 14328
rect 10744 14288 10750 14300
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 900 14232 2360 14260
rect 900 14220 906 14232
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5960 14232 6009 14260
rect 5960 14220 5966 14232
rect 5997 14229 6009 14232
rect 6043 14260 6055 14263
rect 6457 14263 6515 14269
rect 6457 14260 6469 14263
rect 6043 14232 6469 14260
rect 6043 14229 6055 14232
rect 5997 14223 6055 14229
rect 6457 14229 6469 14232
rect 6503 14229 6515 14263
rect 6457 14223 6515 14229
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 12544 14260 12572 14356
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 16132 14328 16160 14359
rect 16942 14356 16948 14408
rect 17000 14356 17006 14408
rect 17052 14396 17080 14436
rect 17310 14424 17316 14476
rect 17368 14424 17374 14476
rect 18322 14424 18328 14476
rect 18380 14424 18386 14476
rect 18969 14467 19027 14473
rect 18969 14433 18981 14467
rect 19015 14433 19027 14467
rect 18969 14427 19027 14433
rect 18874 14396 18880 14408
rect 17052 14368 18880 14396
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 12952 14300 16160 14328
rect 12952 14288 12958 14300
rect 17586 14288 17592 14340
rect 17644 14328 17650 14340
rect 18233 14331 18291 14337
rect 18233 14328 18245 14331
rect 17644 14300 18245 14328
rect 17644 14288 17650 14300
rect 18233 14297 18245 14300
rect 18279 14328 18291 14331
rect 18322 14328 18328 14340
rect 18279 14300 18328 14328
rect 18279 14297 18291 14300
rect 18233 14291 18291 14297
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 18984 14272 19012 14427
rect 10652 14232 12572 14260
rect 10652 14220 10658 14232
rect 12986 14220 12992 14272
rect 13044 14260 13050 14272
rect 15381 14263 15439 14269
rect 15381 14260 15393 14263
rect 13044 14232 15393 14260
rect 13044 14220 13050 14232
rect 15381 14229 15393 14232
rect 15427 14229 15439 14263
rect 15381 14223 15439 14229
rect 16666 14220 16672 14272
rect 16724 14220 16730 14272
rect 18690 14220 18696 14272
rect 18748 14220 18754 14272
rect 18966 14220 18972 14272
rect 19024 14220 19030 14272
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 2130 14016 2136 14068
rect 2188 14016 2194 14068
rect 2590 14016 2596 14068
rect 2648 14056 2654 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2648 14028 2789 14056
rect 2648 14016 2654 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 2777 14019 2835 14025
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 4893 14059 4951 14065
rect 4893 14056 4905 14059
rect 4856 14028 4905 14056
rect 4856 14016 4862 14028
rect 4893 14025 4905 14028
rect 4939 14025 4951 14059
rect 4893 14019 4951 14025
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6052 14028 6377 14056
rect 6052 14016 6058 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9674 14056 9680 14068
rect 9447 14028 9680 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 9824 14028 10548 14056
rect 9824 14016 9830 14028
rect 2148 13988 2176 14016
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 2148 13960 3249 13988
rect 2608 13861 2636 13960
rect 3237 13957 3249 13960
rect 3283 13957 3295 13991
rect 6917 13991 6975 13997
rect 6917 13988 6929 13991
rect 3237 13951 3295 13957
rect 6656 13960 6929 13988
rect 6656 13932 6684 13960
rect 6917 13957 6929 13960
rect 6963 13988 6975 13991
rect 7374 13988 7380 14000
rect 6963 13960 7380 13988
rect 6963 13957 6975 13960
rect 6917 13951 6975 13957
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 7892 13960 9812 13988
rect 7892 13948 7898 13960
rect 3142 13920 3148 13932
rect 2792 13892 3148 13920
rect 2792 13861 2820 13892
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 5534 13920 5540 13932
rect 3252 13892 5540 13920
rect 2593 13855 2651 13861
rect 2593 13821 2605 13855
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2038 13744 2044 13796
rect 2096 13784 2102 13796
rect 3252 13784 3280 13892
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 9784 13920 9812 13960
rect 9953 13923 10011 13929
rect 9953 13920 9965 13923
rect 9784 13892 9965 13920
rect 9953 13889 9965 13892
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 10134 13880 10140 13932
rect 10192 13880 10198 13932
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 4246 13852 4252 13864
rect 3651 13824 4252 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 7006 13852 7012 13864
rect 6227 13824 7012 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7098 13812 7104 13864
rect 7156 13812 7162 13864
rect 7190 13812 7196 13864
rect 7248 13812 7254 13864
rect 7466 13812 7472 13864
rect 7524 13852 7530 13864
rect 9766 13852 9772 13864
rect 7524 13824 9772 13852
rect 7524 13812 7530 13824
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10152 13852 10180 13880
rect 9907 13824 10180 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 10226 13812 10232 13864
rect 10284 13812 10290 13864
rect 10520 13861 10548 14028
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 14369 14059 14427 14065
rect 14369 14056 14381 14059
rect 11020 14028 14381 14056
rect 11020 14016 11026 14028
rect 14369 14025 14381 14028
rect 14415 14025 14427 14059
rect 14369 14019 14427 14025
rect 18874 14016 18880 14068
rect 18932 14016 18938 14068
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 11054 13988 11060 14000
rect 10827 13960 11060 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 15010 13948 15016 14000
rect 15068 13988 15074 14000
rect 15105 13991 15163 13997
rect 15105 13988 15117 13991
rect 15068 13960 15117 13988
rect 15068 13948 15074 13960
rect 15105 13957 15117 13960
rect 15151 13957 15163 13991
rect 15105 13951 15163 13957
rect 15286 13948 15292 14000
rect 15344 13948 15350 14000
rect 14645 13923 14703 13929
rect 10796 13892 12388 13920
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13821 10563 13855
rect 10505 13815 10563 13821
rect 10594 13812 10600 13864
rect 10652 13812 10658 13864
rect 2096 13756 3280 13784
rect 2096 13744 2102 13756
rect 6546 13744 6552 13796
rect 6604 13744 6610 13796
rect 6641 13787 6699 13793
rect 6641 13753 6653 13787
rect 6687 13784 6699 13787
rect 7116 13784 7144 13812
rect 6687 13756 7144 13784
rect 6687 13753 6699 13756
rect 6641 13747 6699 13753
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 10413 13787 10471 13793
rect 9180 13756 9904 13784
rect 9180 13744 9186 13756
rect 6733 13719 6791 13725
rect 6733 13685 6745 13719
rect 6779 13716 6791 13719
rect 6822 13716 6828 13728
rect 6779 13688 6828 13716
rect 6779 13685 6791 13688
rect 6733 13679 6791 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 7009 13719 7067 13725
rect 7009 13685 7021 13719
rect 7055 13716 7067 13719
rect 7098 13716 7104 13728
rect 7055 13688 7104 13716
rect 7055 13685 7067 13688
rect 7009 13679 7067 13685
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 9876 13716 9904 13756
rect 10413 13753 10425 13787
rect 10459 13784 10471 13787
rect 10796 13784 10824 13892
rect 11238 13812 11244 13864
rect 11296 13812 11302 13864
rect 12360 13796 12388 13892
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 15304 13920 15332 13948
rect 14691 13892 15332 13920
rect 16761 13923 16819 13929
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16807 13892 17049 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12618 13852 12624 13864
rect 12483 13824 12624 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12618 13812 12624 13824
rect 12676 13852 12682 13864
rect 12676 13824 13400 13852
rect 12676 13812 12682 13824
rect 13372 13796 13400 13824
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 14516 13824 14565 13852
rect 14516 13812 14522 13824
rect 14553 13821 14565 13824
rect 14599 13852 14611 13855
rect 14918 13852 14924 13864
rect 14599 13824 14924 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 16206 13852 16212 13864
rect 15335 13824 16212 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 16868 13861 16896 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13852 16911 13855
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 16899 13824 17233 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 17221 13821 17233 13824
rect 17267 13852 17279 13855
rect 17586 13852 17592 13864
rect 17267 13824 17592 13852
rect 17267 13821 17279 13824
rect 17221 13815 17279 13821
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 18509 13855 18567 13861
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 18874 13852 18880 13864
rect 18555 13824 18880 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19150 13852 19156 13864
rect 19107 13824 19156 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 10459 13756 10824 13784
rect 11057 13787 11115 13793
rect 10459 13753 10471 13756
rect 10413 13747 10471 13753
rect 11057 13753 11069 13787
rect 11103 13784 11115 13787
rect 11422 13784 11428 13796
rect 11103 13756 11428 13784
rect 11103 13753 11115 13756
rect 11057 13747 11115 13753
rect 10428 13716 10456 13747
rect 11422 13744 11428 13756
rect 11480 13784 11486 13796
rect 12253 13787 12311 13793
rect 12253 13784 12265 13787
rect 11480 13756 12265 13784
rect 11480 13744 11486 13756
rect 12253 13753 12265 13756
rect 12299 13753 12311 13787
rect 12253 13747 12311 13753
rect 9876 13688 10456 13716
rect 10870 13676 10876 13728
rect 10928 13676 10934 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 11388 13688 12081 13716
rect 11388 13676 11394 13688
rect 12069 13685 12081 13688
rect 12115 13685 12127 13719
rect 12268 13716 12296 13747
rect 12342 13744 12348 13796
rect 12400 13744 12406 13796
rect 13354 13744 13360 13796
rect 13412 13744 13418 13796
rect 15105 13787 15163 13793
rect 15105 13753 15117 13787
rect 15151 13784 15163 13787
rect 15194 13784 15200 13796
rect 15151 13756 15200 13784
rect 15151 13753 15163 13756
rect 15105 13747 15163 13753
rect 15194 13744 15200 13756
rect 15252 13784 15258 13796
rect 15562 13784 15568 13796
rect 15252 13756 15568 13784
rect 15252 13744 15258 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 12802 13716 12808 13728
rect 12268 13688 12808 13716
rect 12069 13679 12127 13685
rect 12802 13676 12808 13688
rect 12860 13716 12866 13728
rect 18690 13716 18696 13728
rect 12860 13688 18696 13716
rect 12860 13676 12866 13688
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5994 13521 6000 13524
rect 5461 13515 5519 13521
rect 5461 13512 5473 13515
rect 5040 13484 5473 13512
rect 5040 13472 5046 13484
rect 5461 13481 5473 13484
rect 5507 13481 5519 13515
rect 5461 13475 5519 13481
rect 5981 13515 6000 13521
rect 5981 13481 5993 13515
rect 5981 13475 6000 13481
rect 5994 13472 6000 13475
rect 6052 13472 6058 13524
rect 7466 13512 7472 13524
rect 6104 13484 7472 13512
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 5261 13447 5319 13453
rect 5261 13444 5273 13447
rect 4304 13416 5273 13444
rect 4304 13404 4310 13416
rect 5261 13413 5273 13416
rect 5307 13444 5319 13447
rect 5350 13444 5356 13456
rect 5307 13416 5356 13444
rect 5307 13413 5319 13416
rect 5261 13407 5319 13413
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 6104 13444 6132 13484
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 8665 13515 8723 13521
rect 8665 13481 8677 13515
rect 8711 13512 8723 13515
rect 12342 13512 12348 13524
rect 8711 13484 9444 13512
rect 8711 13481 8723 13484
rect 8665 13475 8723 13481
rect 5552 13416 6132 13444
rect 6181 13447 6239 13453
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 2130 13376 2136 13388
rect 1995 13348 2136 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 2130 13336 2136 13348
rect 2188 13376 2194 13388
rect 3142 13376 3148 13388
rect 2188 13348 3148 13376
rect 2188 13336 2194 13348
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 5166 13336 5172 13388
rect 5224 13336 5230 13388
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2038 13308 2044 13320
rect 1728 13280 2044 13308
rect 1728 13268 1734 13280
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 5552 13308 5580 13416
rect 6181 13413 6193 13447
rect 6227 13444 6239 13447
rect 6730 13444 6736 13456
rect 6227 13416 6736 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 6825 13447 6883 13453
rect 6825 13413 6837 13447
rect 6871 13444 6883 13447
rect 7098 13444 7104 13456
rect 6871 13416 7104 13444
rect 6871 13413 6883 13416
rect 6825 13407 6883 13413
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 7282 13404 7288 13456
rect 7340 13404 7346 13456
rect 8128 13416 8985 13444
rect 6086 13336 6092 13388
rect 6144 13376 6150 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6144 13348 6561 13376
rect 6144 13336 6150 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 6549 13339 6607 13345
rect 4948 13280 5580 13308
rect 4948 13268 4954 13280
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 8128 13308 8156 13416
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8352 13348 8493 13376
rect 8352 13336 8358 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 8662 13336 8668 13388
rect 8720 13336 8726 13388
rect 8957 13385 8985 13416
rect 9122 13404 9128 13456
rect 9180 13404 9186 13456
rect 9416 13444 9444 13484
rect 12084 13484 12348 13512
rect 10686 13444 10692 13456
rect 9416 13416 9536 13444
rect 9508 13388 9536 13416
rect 9784 13416 10692 13444
rect 8838 13379 8896 13385
rect 8838 13376 8850 13379
rect 8772 13348 8850 13376
rect 6880 13280 8156 13308
rect 6880 13268 6886 13280
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8772 13308 8800 13348
rect 8838 13345 8850 13348
rect 8884 13345 8896 13379
rect 8838 13339 8896 13345
rect 8942 13379 9000 13385
rect 8942 13345 8954 13379
rect 8988 13345 9000 13379
rect 8942 13339 9000 13345
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13345 9275 13379
rect 9217 13339 9275 13345
rect 9333 13379 9391 13385
rect 9333 13345 9345 13379
rect 9379 13345 9391 13379
rect 9333 13339 9391 13345
rect 9232 13308 9260 13339
rect 8260 13280 8800 13308
rect 8864 13280 9260 13308
rect 8260 13268 8266 13280
rect 1854 13200 1860 13252
rect 1912 13200 1918 13252
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 5629 13243 5687 13249
rect 4580 13212 5580 13240
rect 4580 13200 4586 13212
rect 1762 13132 1768 13184
rect 1820 13132 1826 13184
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 3568 13144 4261 13172
rect 3568 13132 3574 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4249 13135 4307 13141
rect 4982 13132 4988 13184
rect 5040 13132 5046 13184
rect 5442 13132 5448 13184
rect 5500 13132 5506 13184
rect 5552 13172 5580 13212
rect 5629 13209 5641 13243
rect 5675 13240 5687 13243
rect 5675 13212 6040 13240
rect 5675 13209 5687 13212
rect 5629 13203 5687 13209
rect 6012 13181 6040 13212
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5552 13144 5825 13172
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 5813 13135 5871 13141
rect 5997 13175 6055 13181
rect 5997 13141 6009 13175
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 8297 13175 8355 13181
rect 8297 13172 8309 13175
rect 8168 13144 8309 13172
rect 8168 13132 8174 13144
rect 8297 13141 8309 13144
rect 8343 13141 8355 13175
rect 8864 13172 8892 13280
rect 8938 13200 8944 13252
rect 8996 13240 9002 13252
rect 9348 13240 9376 13339
rect 9490 13336 9496 13388
rect 9548 13380 9554 13388
rect 9784 13385 9812 13416
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 12084 13453 12112 13484
rect 12342 13472 12348 13484
rect 12400 13512 12406 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 12400 13484 13553 13512
rect 12400 13472 12406 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 13541 13475 13599 13481
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 14090 13512 14096 13524
rect 13771 13484 14096 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 14090 13472 14096 13484
rect 14148 13512 14154 13524
rect 14148 13484 15056 13512
rect 14148 13472 14154 13484
rect 12069 13447 12127 13453
rect 12069 13413 12081 13447
rect 12115 13413 12127 13447
rect 12069 13407 12127 13413
rect 14277 13447 14335 13453
rect 14277 13413 14289 13447
rect 14323 13444 14335 13447
rect 14323 13416 14964 13444
rect 14323 13413 14335 13416
rect 14277 13407 14335 13413
rect 9585 13380 9643 13385
rect 9548 13379 9643 13380
rect 9548 13352 9597 13379
rect 9548 13336 9554 13352
rect 9585 13345 9597 13352
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10870 13376 10876 13388
rect 10183 13348 10876 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11146 13336 11152 13388
rect 11204 13336 11210 13388
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11425 13379 11483 13385
rect 11296 13348 11341 13376
rect 11296 13336 11302 13348
rect 11425 13345 11437 13379
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 10042 13268 10048 13320
rect 10100 13268 10106 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10502 13308 10508 13320
rect 10284 13280 10508 13308
rect 10284 13268 10290 13280
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 11440 13308 11468 13339
rect 11514 13336 11520 13388
rect 11572 13336 11578 13388
rect 11698 13385 11704 13388
rect 11655 13379 11704 13385
rect 11655 13345 11667 13379
rect 11701 13345 11704 13379
rect 11655 13339 11704 13345
rect 11698 13336 11704 13339
rect 11756 13336 11762 13388
rect 11882 13336 11888 13388
rect 11940 13336 11946 13388
rect 12158 13336 12164 13388
rect 12216 13336 12222 13388
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13376 12311 13379
rect 12526 13376 12532 13388
rect 12299 13348 12532 13376
rect 12299 13345 12311 13348
rect 12253 13339 12311 13345
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 12894 13336 12900 13388
rect 12952 13336 12958 13388
rect 12986 13336 12992 13388
rect 13044 13336 13050 13388
rect 13078 13336 13084 13388
rect 13136 13336 13142 13388
rect 13170 13336 13176 13388
rect 13228 13385 13234 13388
rect 13228 13379 13257 13385
rect 13245 13345 13257 13379
rect 13228 13339 13257 13345
rect 13228 13336 13234 13339
rect 13354 13336 13360 13388
rect 13412 13336 13418 13388
rect 14458 13336 14464 13388
rect 14516 13336 14522 13388
rect 13188 13308 13216 13336
rect 11440 13280 13216 13308
rect 13817 13311 13875 13317
rect 8996 13212 9376 13240
rect 8996 13200 9002 13212
rect 9858 13200 9864 13252
rect 9916 13240 9922 13252
rect 11440 13240 11468 13280
rect 13817 13277 13829 13311
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 9916 13212 11468 13240
rect 9916 13200 9922 13212
rect 13832 13184 13860 13271
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 14476 13240 14504 13336
rect 14936 13308 14964 13416
rect 15028 13388 15056 13484
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 17957 13515 18015 13521
rect 17957 13512 17969 13515
rect 17552 13484 17969 13512
rect 17552 13472 17558 13484
rect 17957 13481 17969 13484
rect 18003 13481 18015 13515
rect 17957 13475 18015 13481
rect 16206 13444 16212 13456
rect 16132 13416 16212 13444
rect 15010 13336 15016 13388
rect 15068 13336 15074 13388
rect 15286 13376 15292 13388
rect 15166 13348 15292 13376
rect 15166 13308 15194 13348
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15562 13336 15568 13388
rect 15620 13336 15626 13388
rect 16132 13385 16160 13416
rect 16206 13404 16212 13416
rect 16264 13444 16270 13456
rect 17512 13444 17540 13472
rect 16264 13416 17540 13444
rect 16264 13404 16270 13416
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 15672 13308 15700 13339
rect 17586 13336 17592 13388
rect 17644 13336 17650 13388
rect 18230 13336 18236 13388
rect 18288 13336 18294 13388
rect 14936 13280 15700 13308
rect 17604 13249 17632 13336
rect 14332 13212 14504 13240
rect 17589 13243 17647 13249
rect 14332 13200 14338 13212
rect 17589 13209 17601 13243
rect 17635 13240 17647 13243
rect 17862 13240 17868 13252
rect 17635 13212 17868 13240
rect 17635 13209 17647 13212
rect 17589 13203 17647 13209
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 9306 13172 9312 13184
rect 8864 13144 9312 13172
rect 8297 13135 8355 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9493 13175 9551 13181
rect 9493 13141 9505 13175
rect 9539 13172 9551 13175
rect 10962 13172 10968 13184
rect 9539 13144 10968 13172
rect 9539 13141 9551 13144
rect 9493 13135 9551 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 11974 13172 11980 13184
rect 11839 13144 11980 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12437 13175 12495 13181
rect 12437 13141 12449 13175
rect 12483 13172 12495 13175
rect 12526 13172 12532 13184
rect 12483 13144 12532 13172
rect 12483 13141 12495 13144
rect 12437 13135 12495 13141
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 13814 13132 13820 13184
rect 13872 13132 13878 13184
rect 14550 13132 14556 13184
rect 14608 13132 14614 13184
rect 18598 13132 18604 13184
rect 18656 13132 18662 13184
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 2869 12971 2927 12977
rect 2869 12968 2881 12971
rect 2648 12940 2881 12968
rect 2648 12928 2654 12940
rect 2869 12937 2881 12940
rect 2915 12968 2927 12971
rect 4798 12968 4804 12980
rect 2915 12940 4108 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 3142 12860 3148 12912
rect 3200 12900 3206 12912
rect 3200 12872 3648 12900
rect 3200 12860 3206 12872
rect 1121 12835 1179 12841
rect 1121 12801 1133 12835
rect 1167 12832 1179 12835
rect 1762 12832 1768 12844
rect 1167 12804 1768 12832
rect 1167 12801 1179 12804
rect 1121 12795 1179 12801
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 842 12724 848 12776
rect 900 12724 906 12776
rect 3510 12724 3516 12776
rect 3568 12724 3574 12776
rect 3620 12773 3648 12872
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3694 12724 3700 12776
rect 3752 12724 3758 12776
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 3970 12764 3976 12776
rect 3927 12736 3976 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 2498 12696 2504 12708
rect 2346 12668 2504 12696
rect 2498 12656 2504 12668
rect 2556 12656 2562 12708
rect 2682 12656 2688 12708
rect 2740 12656 2746 12708
rect 2901 12699 2959 12705
rect 2901 12665 2913 12699
rect 2947 12696 2959 12699
rect 2947 12668 3832 12696
rect 2947 12665 2959 12668
rect 2901 12659 2959 12665
rect 3804 12640 3832 12668
rect 3050 12588 3056 12640
rect 3108 12588 3114 12640
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 3786 12588 3792 12640
rect 3844 12588 3850 12640
rect 4080 12628 4108 12940
rect 4356 12940 4804 12968
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4356 12841 4384 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 5224 12940 6193 12968
rect 5224 12928 5230 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 7190 12928 7196 12980
rect 7248 12928 7254 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 10229 12971 10287 12977
rect 8720 12940 9674 12968
rect 8720 12928 8726 12940
rect 8110 12900 8116 12912
rect 7668 12872 8116 12900
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4212 12804 4353 12832
rect 4212 12792 4218 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4982 12832 4988 12844
rect 4663 12804 4988 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 6089 12835 6147 12841
rect 5316 12804 5948 12832
rect 5316 12792 5322 12804
rect 4338 12656 4344 12708
rect 4396 12696 4402 12708
rect 5920 12696 5948 12804
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 6135 12804 6653 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 6656 12764 6684 12795
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 7668 12841 7696 12872
rect 8110 12860 8116 12872
rect 8168 12900 8174 12912
rect 9398 12900 9404 12912
rect 8168 12872 9404 12900
rect 8168 12860 8174 12872
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 9490 12860 9496 12912
rect 9548 12860 9554 12912
rect 7653 12835 7711 12841
rect 6880 12804 7604 12832
rect 6880 12792 6886 12804
rect 7190 12764 7196 12776
rect 6656 12736 7196 12764
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7576 12764 7604 12804
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 7834 12792 7840 12844
rect 7892 12792 7898 12844
rect 8496 12804 8708 12832
rect 7852 12764 7880 12792
rect 8496 12776 8524 12804
rect 7576 12736 7880 12764
rect 8478 12724 8484 12776
rect 8536 12724 8542 12776
rect 8570 12724 8576 12776
rect 8628 12724 8634 12776
rect 8680 12773 8708 12804
rect 8846 12792 8852 12844
rect 8904 12792 8910 12844
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9508 12832 9536 12860
rect 9324 12804 9536 12832
rect 9646 12832 9674 12940
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 10318 12968 10324 12980
rect 10275 12940 10324 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11330 12968 11336 12980
rect 10520 12940 11336 12968
rect 9766 12832 9772 12844
rect 9646 12804 9772 12832
rect 8666 12767 8724 12773
rect 8666 12733 8678 12767
rect 8712 12733 8724 12767
rect 8864 12764 8892 12792
rect 8666 12727 8724 12733
rect 8772 12736 8892 12764
rect 8956 12764 8984 12792
rect 9324 12776 9352 12804
rect 9766 12792 9772 12804
rect 9824 12832 9830 12844
rect 10042 12832 10048 12844
rect 9824 12804 10048 12832
rect 9824 12792 9830 12804
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 9038 12767 9096 12773
rect 9038 12764 9050 12767
rect 8956 12736 9050 12764
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 4396 12668 5106 12696
rect 5920 12668 7573 12696
rect 4396 12656 4402 12668
rect 7561 12665 7573 12668
rect 7607 12696 7619 12699
rect 8772 12696 8800 12736
rect 9038 12733 9050 12736
rect 9084 12733 9096 12767
rect 9038 12727 9096 12733
rect 9214 12724 9220 12776
rect 9272 12724 9278 12776
rect 9306 12724 9312 12776
rect 9364 12724 9370 12776
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9456 12736 9505 12764
rect 9456 12724 9462 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 9909 12767 9967 12773
rect 9909 12733 9921 12767
rect 9955 12764 9967 12767
rect 10520 12764 10548 12940
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 11606 12928 11612 12980
rect 11664 12928 11670 12980
rect 12526 12928 12532 12980
rect 12584 12928 12590 12980
rect 12621 12971 12679 12977
rect 12621 12937 12633 12971
rect 12667 12968 12679 12971
rect 12710 12968 12716 12980
rect 12667 12940 12716 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 10686 12860 10692 12912
rect 10744 12860 10750 12912
rect 10870 12860 10876 12912
rect 10928 12900 10934 12912
rect 11149 12903 11207 12909
rect 10928 12872 11008 12900
rect 10928 12860 10934 12872
rect 9955 12736 10548 12764
rect 10597 12767 10655 12773
rect 9955 12733 9967 12736
rect 9909 12727 9967 12733
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 10704 12764 10732 12860
rect 10778 12792 10784 12844
rect 10836 12792 10842 12844
rect 10643 12736 10732 12764
rect 10796 12764 10824 12792
rect 10980 12773 11008 12872
rect 11149 12869 11161 12903
rect 11195 12869 11207 12903
rect 11149 12863 11207 12869
rect 11164 12832 11192 12863
rect 12342 12860 12348 12912
rect 12400 12900 12406 12912
rect 12986 12900 12992 12912
rect 12400 12872 12992 12900
rect 12400 12860 12406 12872
rect 12986 12860 12992 12872
rect 13044 12860 13050 12912
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 15562 12900 15568 12912
rect 13872 12872 15568 12900
rect 13872 12860 13878 12872
rect 14090 12841 14096 12844
rect 11425 12835 11483 12841
rect 11425 12832 11437 12835
rect 11164 12804 11437 12832
rect 11425 12801 11437 12804
rect 11471 12801 11483 12835
rect 11425 12795 11483 12801
rect 14068 12835 14096 12841
rect 14068 12801 14080 12835
rect 14068 12795 14096 12801
rect 14090 12792 14096 12795
rect 14148 12792 14154 12844
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14274 12832 14280 12844
rect 14231 12804 14280 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14568 12841 14596 12872
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 15013 12835 15071 12841
rect 15013 12801 15025 12835
rect 15059 12832 15071 12835
rect 15059 12804 15148 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 15120 12776 15148 12804
rect 16206 12792 16212 12844
rect 16264 12792 16270 12844
rect 17773 12835 17831 12841
rect 17773 12801 17785 12835
rect 17819 12832 17831 12835
rect 17819 12804 17908 12832
rect 17819 12801 17831 12804
rect 17773 12795 17831 12801
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10796 12736 10885 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 7607 12668 8800 12696
rect 8849 12699 8907 12705
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 8849 12665 8861 12699
rect 8895 12665 8907 12699
rect 8849 12659 8907 12665
rect 8941 12699 8999 12705
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 9232 12696 9260 12724
rect 8987 12668 9260 12696
rect 9508 12696 9536 12727
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11333 12767 11391 12773
rect 11333 12764 11345 12767
rect 11112 12736 11345 12764
rect 11112 12724 11118 12736
rect 11333 12733 11345 12736
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 11514 12724 11520 12776
rect 11572 12764 11578 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11572 12736 11621 12764
rect 11572 12724 11578 12736
rect 11609 12733 11621 12736
rect 11655 12764 11667 12767
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 11655 12736 12725 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 12802 12724 12808 12776
rect 12860 12724 12866 12776
rect 12986 12724 12992 12776
rect 13044 12724 13050 12776
rect 15102 12724 15108 12776
rect 15160 12724 15166 12776
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16482 12764 16488 12776
rect 16347 12736 16488 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 17880 12773 17908 12804
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18656 12804 19073 12832
rect 18656 12792 18662 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12733 17923 12767
rect 17865 12727 17923 12733
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 9508 12668 10548 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 5258 12628 5264 12640
rect 4080 12600 5264 12628
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 5408 12600 6561 12628
rect 5408 12588 5414 12600
rect 6549 12597 6561 12600
rect 6595 12628 6607 12631
rect 7834 12628 7840 12640
rect 6595 12600 7840 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8864 12628 8892 12659
rect 10520 12640 10548 12668
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 10836 12668 13216 12696
rect 10836 12656 10842 12668
rect 9122 12628 9128 12640
rect 8864 12600 9128 12628
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9217 12631 9275 12637
rect 9217 12597 9229 12631
rect 9263 12628 9275 12631
rect 9490 12628 9496 12640
rect 9263 12600 9496 12628
rect 9263 12597 9275 12600
rect 9217 12591 9275 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 9766 12628 9772 12640
rect 9640 12600 9772 12628
rect 9640 12588 9646 12600
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 10502 12588 10508 12640
rect 10560 12588 10566 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 12066 12628 12072 12640
rect 11839 12600 12072 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12526 12628 12532 12640
rect 12299 12600 12532 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 13188 12628 13216 12668
rect 13538 12656 13544 12708
rect 13596 12656 13602 12708
rect 13725 12699 13783 12705
rect 13725 12665 13737 12699
rect 13771 12696 13783 12699
rect 13771 12668 14320 12696
rect 13771 12665 13783 12668
rect 13725 12659 13783 12665
rect 14292 12637 14320 12668
rect 17880 12640 17908 12727
rect 13909 12631 13967 12637
rect 13909 12628 13921 12631
rect 13188 12600 13921 12628
rect 13909 12597 13921 12600
rect 13955 12597 13967 12631
rect 13909 12591 13967 12597
rect 14277 12631 14335 12637
rect 14277 12597 14289 12631
rect 14323 12628 14335 12631
rect 15286 12628 15292 12640
rect 14323 12600 15292 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 17862 12588 17868 12640
rect 17920 12628 17926 12640
rect 18708 12637 18736 12727
rect 18693 12631 18751 12637
rect 18693 12628 18705 12631
rect 17920 12600 18705 12628
rect 17920 12588 17926 12600
rect 18693 12597 18705 12600
rect 18739 12597 18751 12631
rect 18693 12591 18751 12597
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 3694 12424 3700 12436
rect 1780 12396 3004 12424
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 1780 12297 1808 12396
rect 2516 12365 2544 12396
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2480 12359 2544 12365
rect 1903 12328 2452 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 1728 12260 1777 12288
rect 1728 12248 1734 12260
rect 1765 12257 1777 12260
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12288 2099 12291
rect 2424 12288 2452 12328
rect 2480 12325 2492 12359
rect 2526 12328 2544 12359
rect 2682 12356 2688 12368
rect 2608 12328 2688 12356
rect 2526 12325 2538 12328
rect 2480 12319 2538 12325
rect 2608 12288 2636 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 2976 12297 3004 12396
rect 3068 12396 3700 12424
rect 2087 12260 2360 12288
rect 2087 12257 2099 12260
rect 2041 12251 2099 12257
rect 2130 12180 2136 12232
rect 2188 12180 2194 12232
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 2041 12155 2099 12161
rect 2041 12152 2053 12155
rect 1912 12124 2053 12152
rect 1912 12112 1918 12124
rect 2041 12121 2053 12124
rect 2087 12121 2099 12155
rect 2041 12115 2099 12121
rect 2148 12084 2176 12180
rect 2332 12152 2360 12260
rect 2424 12260 2636 12288
rect 2777 12291 2835 12297
rect 2424 12232 2452 12260
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 2406 12180 2412 12232
rect 2464 12180 2470 12232
rect 2792 12152 2820 12251
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3068 12220 3096 12396
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 3786 12384 3792 12436
rect 3844 12424 3850 12436
rect 4890 12424 4896 12436
rect 3844 12396 4896 12424
rect 3844 12384 3850 12396
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 8260 12396 8401 12424
rect 8260 12384 8266 12396
rect 8389 12393 8401 12396
rect 8435 12393 8447 12427
rect 10594 12424 10600 12436
rect 8389 12387 8447 12393
rect 8496 12396 10600 12424
rect 3418 12316 3424 12368
rect 3476 12316 3482 12368
rect 7377 12359 7435 12365
rect 7377 12325 7389 12359
rect 7423 12356 7435 12359
rect 7423 12328 7696 12356
rect 7423 12325 7435 12328
rect 7377 12319 7435 12325
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4488 12260 4554 12288
rect 4488 12248 4494 12260
rect 6454 12248 6460 12300
rect 6512 12248 6518 12300
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 6696 12260 7205 12288
rect 6696 12248 6702 12260
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7668 12288 7696 12328
rect 7668 12260 7788 12288
rect 7561 12251 7619 12257
rect 2915 12192 3096 12220
rect 3145 12223 3203 12229
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3145 12189 3157 12223
rect 3191 12189 3203 12223
rect 7576 12220 7604 12251
rect 7760 12220 7788 12260
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 8018 12248 8024 12300
rect 8076 12248 8082 12300
rect 8110 12248 8116 12300
rect 8168 12248 8174 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12257 8263 12291
rect 8205 12251 8263 12257
rect 8036 12220 8064 12248
rect 7576 12192 7696 12220
rect 7760 12192 8064 12220
rect 8220 12220 8248 12251
rect 8496 12220 8524 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11664 12396 11805 12424
rect 11664 12384 11670 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 11961 12427 12019 12433
rect 11961 12393 11973 12427
rect 12007 12424 12019 12427
rect 12618 12424 12624 12436
rect 12007 12396 12624 12424
rect 12007 12393 12019 12396
rect 11961 12387 12019 12393
rect 12618 12384 12624 12396
rect 12676 12424 12682 12436
rect 12894 12424 12900 12436
rect 12676 12396 12900 12424
rect 12676 12384 12682 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13170 12384 13176 12436
rect 13228 12384 13234 12436
rect 13541 12427 13599 12433
rect 13541 12424 13553 12427
rect 13280 12396 13553 12424
rect 9030 12316 9036 12368
rect 9088 12316 9094 12368
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 11054 12356 11060 12368
rect 9180 12328 11060 12356
rect 9180 12316 9186 12328
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 12158 12356 12164 12368
rect 11296 12328 12164 12356
rect 11296 12316 11302 12328
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 13280 12356 13308 12396
rect 13541 12393 13553 12396
rect 13587 12424 13599 12427
rect 15194 12424 15200 12436
rect 13587 12396 15200 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 15194 12384 15200 12396
rect 15252 12424 15258 12436
rect 16666 12424 16672 12436
rect 15252 12396 16672 12424
rect 15252 12384 15258 12396
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 12912 12328 13308 12356
rect 13449 12359 13507 12365
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9272 12260 9505 12288
rect 9272 12248 9278 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9692 12220 9720 12251
rect 10042 12248 10048 12300
rect 10100 12248 10106 12300
rect 11422 12248 11428 12300
rect 11480 12248 11486 12300
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 11790 12288 11796 12300
rect 11747 12260 11796 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 12342 12288 12348 12300
rect 11900 12260 12348 12288
rect 8220 12192 8524 12220
rect 9140 12192 9720 12220
rect 9953 12223 10011 12229
rect 3145 12183 3203 12189
rect 3050 12152 3056 12164
rect 2332 12124 2544 12152
rect 2792 12124 3056 12152
rect 2516 12093 2544 12124
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 2148 12056 2329 12084
rect 2317 12053 2329 12056
rect 2363 12053 2375 12087
rect 2317 12047 2375 12053
rect 2501 12087 2559 12093
rect 2501 12053 2513 12087
rect 2547 12084 2559 12087
rect 2590 12084 2596 12096
rect 2547 12056 2596 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 3160 12084 3188 12183
rect 7668 12152 7696 12192
rect 8220 12152 8248 12192
rect 9140 12164 9168 12192
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 7668 12124 8248 12152
rect 9122 12112 9128 12164
rect 9180 12112 9186 12164
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9674 12152 9680 12164
rect 9364 12124 9680 12152
rect 9364 12112 9370 12124
rect 9674 12112 9680 12124
rect 9732 12152 9738 12164
rect 9968 12152 9996 12183
rect 9732 12124 9996 12152
rect 9732 12112 9738 12124
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 11425 12155 11483 12161
rect 11425 12152 11437 12155
rect 11112 12124 11437 12152
rect 11112 12112 11118 12124
rect 11425 12121 11437 12124
rect 11471 12121 11483 12155
rect 11425 12115 11483 12121
rect 4154 12084 4160 12096
rect 3160 12056 4160 12084
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 6273 12087 6331 12093
rect 6273 12084 6285 12087
rect 6236 12056 6285 12084
rect 6236 12044 6242 12056
rect 6273 12053 6285 12056
rect 6319 12053 6331 12087
rect 6273 12047 6331 12053
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 9214 12084 9220 12096
rect 7791 12056 9220 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10778 12084 10784 12096
rect 10376 12056 10784 12084
rect 10376 12044 10382 12056
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 11900 12084 11928 12260
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 12912 12288 12940 12328
rect 13449 12325 13461 12359
rect 13495 12356 13507 12359
rect 13814 12356 13820 12368
rect 13495 12328 13820 12356
rect 13495 12325 13507 12328
rect 13449 12319 13507 12325
rect 12483 12260 12572 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12250 12112 12256 12164
rect 12308 12112 12314 12164
rect 12544 12093 12572 12260
rect 12820 12260 12940 12288
rect 12989 12291 13047 12297
rect 12820 12229 12848 12260
rect 12989 12257 13001 12291
rect 13035 12288 13047 12291
rect 13464 12288 13492 12319
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 13035 12260 13492 12288
rect 13035 12257 13047 12260
rect 12989 12251 13047 12257
rect 15102 12248 15108 12300
rect 15160 12288 15166 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15160 12260 15485 12288
rect 15160 12248 15166 12260
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 16393 12291 16451 12297
rect 16393 12288 16405 12291
rect 15620 12260 16405 12288
rect 15620 12248 15626 12260
rect 16393 12257 16405 12260
rect 16439 12257 16451 12291
rect 16393 12251 16451 12257
rect 17862 12248 17868 12300
rect 17920 12248 17926 12300
rect 13354 12229 13360 12232
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13332 12223 13360 12229
rect 13332 12189 13344 12223
rect 13332 12183 13360 12189
rect 12728 12152 12756 12183
rect 12912 12152 12940 12183
rect 13354 12180 13360 12183
rect 13412 12180 13418 12232
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12220 13875 12223
rect 13998 12220 14004 12232
rect 13863 12192 14004 12220
rect 13863 12189 13875 12192
rect 13817 12183 13875 12189
rect 13832 12152 13860 12183
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 15286 12220 15292 12232
rect 14415 12192 15292 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 12728 12124 12848 12152
rect 12912 12124 13860 12152
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11900 12056 11989 12084
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12710 12084 12716 12096
rect 12575 12056 12716 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12820 12084 12848 12124
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 15396 12152 15424 12183
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 18874 12220 18880 12232
rect 16540 12192 18880 12220
rect 16540 12180 16546 12192
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 15160 12124 15424 12152
rect 17773 12155 17831 12161
rect 15160 12112 15166 12124
rect 17773 12121 17785 12155
rect 17819 12152 17831 12155
rect 17862 12152 17868 12164
rect 17819 12124 17868 12152
rect 17819 12121 17831 12124
rect 17773 12115 17831 12121
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 13354 12084 13360 12096
rect 12820 12056 13360 12084
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 16209 12087 16267 12093
rect 16209 12053 16221 12087
rect 16255 12084 16267 12087
rect 16298 12084 16304 12096
rect 16255 12056 16304 12084
rect 16255 12053 16267 12056
rect 16209 12047 16267 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 4709 11883 4767 11889
rect 4709 11849 4721 11883
rect 4755 11880 4767 11883
rect 4798 11880 4804 11892
rect 4755 11852 4804 11880
rect 4755 11849 4767 11852
rect 4709 11843 4767 11849
rect 1486 11772 1492 11824
rect 1544 11772 1550 11824
rect 2961 11815 3019 11821
rect 2961 11781 2973 11815
rect 3007 11812 3019 11815
rect 3326 11812 3332 11824
rect 3007 11784 3332 11812
rect 3007 11781 3019 11784
rect 2961 11775 3019 11781
rect 3326 11772 3332 11784
rect 3384 11772 3390 11824
rect 1688 11716 2452 11744
rect 1489 11679 1547 11685
rect 1489 11645 1501 11679
rect 1535 11676 1547 11679
rect 1578 11676 1584 11688
rect 1535 11648 1584 11676
rect 1535 11645 1547 11648
rect 1489 11639 1547 11645
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 1688 11685 1716 11716
rect 2424 11688 2452 11716
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11645 1731 11679
rect 1673 11639 1731 11645
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 1811 11648 1845 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 1780 11608 1808 11639
rect 2406 11636 2412 11688
rect 2464 11636 2470 11688
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 3234 11676 3240 11688
rect 2731 11648 3240 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11676 4491 11679
rect 4724 11676 4752 11843
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 10045 11883 10103 11889
rect 7616 11852 9904 11880
rect 7616 11840 7622 11852
rect 9876 11812 9904 11852
rect 10045 11849 10057 11883
rect 10091 11880 10103 11883
rect 10410 11880 10416 11892
rect 10091 11852 10416 11880
rect 10091 11849 10103 11852
rect 10045 11843 10103 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 9876 11784 10088 11812
rect 10060 11756 10088 11784
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 13078 11812 13084 11824
rect 12492 11784 13084 11812
rect 12492 11772 12498 11784
rect 13078 11772 13084 11784
rect 13136 11772 13142 11824
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11744 6147 11747
rect 6178 11744 6184 11756
rect 6135 11716 6184 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 9398 11704 9404 11756
rect 9456 11704 9462 11756
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 10042 11704 10048 11756
rect 10100 11704 10106 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14200 11716 14289 11744
rect 4479 11648 4752 11676
rect 4479 11645 4491 11648
rect 4433 11639 4491 11645
rect 4890 11636 4896 11688
rect 4948 11636 4954 11688
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 5040 11648 5181 11676
rect 5040 11636 5046 11648
rect 5169 11645 5181 11648
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 8662 11636 8668 11688
rect 8720 11636 8726 11688
rect 9306 11636 9312 11688
rect 9364 11636 9370 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 11054 11676 11060 11688
rect 9723 11648 11060 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 2777 11611 2835 11617
rect 2777 11608 2789 11611
rect 1688 11580 2789 11608
rect 1688 11552 1716 11580
rect 2777 11577 2789 11580
rect 2823 11577 2835 11611
rect 2777 11571 2835 11577
rect 2961 11611 3019 11617
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 4614 11608 4620 11620
rect 3007 11580 4620 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 1670 11500 1676 11552
rect 1728 11500 1734 11552
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 2976 11540 3004 11571
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 6546 11568 6552 11620
rect 6604 11568 6610 11620
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 8938 11608 8944 11620
rect 8527 11580 8944 11608
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 9692 11608 9720 11639
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11238 11636 11244 11688
rect 11296 11636 11302 11688
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11480 11648 11621 11676
rect 11480 11636 11486 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11756 11648 11805 11676
rect 11756 11636 11762 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 12802 11636 12808 11688
rect 12860 11676 12866 11688
rect 13538 11676 13544 11688
rect 12860 11648 13544 11676
rect 12860 11636 12866 11648
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 14200 11685 14228 11716
rect 14277 11713 14289 11716
rect 14323 11744 14335 11747
rect 15102 11744 15108 11756
rect 14323 11716 15108 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 15102 11704 15108 11716
rect 15160 11744 15166 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 15160 11716 16957 11744
rect 15160 11704 15166 11716
rect 16945 11713 16957 11716
rect 16991 11744 17003 11747
rect 16991 11716 17908 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15344 11648 15393 11676
rect 15344 11636 15350 11648
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 15427 11648 15485 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15473 11645 15485 11648
rect 15519 11676 15531 11679
rect 16482 11676 16488 11688
rect 15519 11648 16488 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 17052 11685 17080 11716
rect 17880 11688 17908 11716
rect 17037 11679 17095 11685
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 17083 11648 17117 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 17310 11636 17316 11688
rect 17368 11636 17374 11688
rect 17862 11636 17868 11688
rect 17920 11636 17926 11688
rect 19058 11636 19064 11688
rect 19116 11636 19122 11688
rect 11514 11608 11520 11620
rect 9140 11580 9720 11608
rect 9784 11580 11520 11608
rect 9140 11552 9168 11580
rect 2648 11512 3004 11540
rect 4341 11543 4399 11549
rect 2648 11500 2654 11512
rect 4341 11509 4353 11543
rect 4387 11540 4399 11543
rect 4430 11540 4436 11552
rect 4387 11512 4436 11540
rect 4387 11509 4399 11512
rect 4341 11503 4399 11509
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4856 11512 4997 11540
rect 4856 11500 4862 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 8110 11540 8116 11552
rect 5500 11512 8116 11540
rect 5500 11500 5506 11512
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8846 11500 8852 11552
rect 8904 11500 8910 11552
rect 9122 11500 9128 11552
rect 9180 11500 9186 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9784 11540 9812 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 12253 11611 12311 11617
rect 12253 11577 12265 11611
rect 12299 11608 12311 11611
rect 15102 11608 15108 11620
rect 12299 11580 15108 11608
rect 12299 11577 12311 11580
rect 12253 11571 12311 11577
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 17126 11568 17132 11620
rect 17184 11568 17190 11620
rect 9456 11512 9812 11540
rect 9456 11500 9462 11512
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 12618 11540 12624 11552
rect 10836 11512 12624 11540
rect 10836 11500 10842 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 14182 11540 14188 11552
rect 13412 11512 14188 11540
rect 13412 11500 13418 11512
rect 14182 11500 14188 11512
rect 14240 11540 14246 11552
rect 15010 11540 15016 11552
rect 14240 11512 15016 11540
rect 14240 11500 14246 11512
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 17368 11512 18889 11540
rect 17368 11500 17374 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 4154 11336 4160 11348
rect 860 11308 4160 11336
rect 860 11212 888 11308
rect 2498 11268 2504 11280
rect 2346 11240 2504 11268
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 842 11160 848 11212
rect 900 11160 906 11212
rect 2884 11209 2912 11308
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4893 11339 4951 11345
rect 4893 11305 4905 11339
rect 4939 11336 4951 11339
rect 4982 11336 4988 11348
rect 4939 11308 4988 11336
rect 4939 11305 4951 11308
rect 4893 11299 4951 11305
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5442 11336 5448 11348
rect 5307 11308 5448 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6454 11296 6460 11348
rect 6512 11296 6518 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7558 11336 7564 11348
rect 6963 11308 7564 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 8297 11339 8355 11345
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 8662 11336 8668 11348
rect 8343 11308 8668 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 8846 11296 8852 11348
rect 8904 11296 8910 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9398 11336 9404 11348
rect 9088 11308 9404 11336
rect 9088 11296 9094 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 9732 11308 9904 11336
rect 9732 11296 9738 11308
rect 4430 11268 4436 11280
rect 4370 11240 4436 11268
rect 4430 11228 4436 11240
rect 4488 11268 4494 11280
rect 6546 11268 6552 11280
rect 4488 11240 6552 11268
rect 4488 11228 4494 11240
rect 6546 11228 6552 11240
rect 6604 11228 6610 11280
rect 6825 11271 6883 11277
rect 6825 11237 6837 11271
rect 6871 11268 6883 11271
rect 7374 11268 7380 11280
rect 6871 11240 7380 11268
rect 6871 11237 6883 11240
rect 6825 11231 6883 11237
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11169 2927 11203
rect 2869 11163 2927 11169
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5994 11200 6000 11212
rect 5399 11172 6000 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 1118 11092 1124 11144
rect 1176 11092 1182 11144
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11132 5595 11135
rect 6822 11132 6828 11144
rect 5583 11104 6828 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6880 11104 7021 11132
rect 6880 11092 6886 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 7116 11064 7144 11240
rect 7374 11228 7380 11240
rect 7432 11228 7438 11280
rect 8036 11240 8248 11268
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 8036 11200 8064 11240
rect 8220 11209 8248 11240
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 8757 11271 8815 11277
rect 8757 11268 8769 11271
rect 8444 11240 8769 11268
rect 8444 11228 8450 11240
rect 8757 11237 8769 11240
rect 8803 11237 8815 11271
rect 8757 11231 8815 11237
rect 7248 11172 8064 11200
rect 8113 11203 8171 11209
rect 7248 11160 7254 11172
rect 4672 11036 7144 11064
rect 4672 11024 4678 11036
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 2593 10999 2651 11005
rect 2593 10996 2605 10999
rect 2464 10968 2605 10996
rect 2464 10956 2470 10968
rect 2593 10965 2605 10968
rect 2639 10996 2651 10999
rect 5442 10996 5448 11008
rect 2639 10968 5448 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 7944 10996 7972 11172
rect 8113 11169 8125 11203
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8128 11132 8156 11163
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8352 11172 8493 11200
rect 8352 11160 8358 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 8864 11200 8892 11296
rect 9876 11209 9904 11308
rect 10226 11296 10232 11348
rect 10284 11296 10290 11348
rect 11054 11296 11060 11348
rect 11112 11296 11118 11348
rect 12434 11336 12440 11348
rect 12406 11296 12440 11336
rect 12492 11296 12498 11348
rect 17402 11336 17408 11348
rect 12636 11308 17408 11336
rect 10244 11268 10272 11296
rect 10321 11271 10379 11277
rect 10321 11268 10333 11271
rect 10244 11240 10333 11268
rect 10321 11237 10333 11240
rect 10367 11237 10379 11271
rect 10321 11231 10379 11237
rect 10410 11228 10416 11280
rect 10468 11268 10474 11280
rect 10686 11268 10692 11280
rect 10468 11240 10692 11268
rect 10468 11228 10474 11240
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 10778 11228 10784 11280
rect 10836 11228 10842 11280
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 8864 11172 9413 11200
rect 8481 11163 8539 11169
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 9122 11132 9128 11144
rect 8128 11104 9128 11132
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9784 11132 9812 11163
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10226 11209 10232 11212
rect 10203 11203 10232 11209
rect 10203 11169 10215 11203
rect 10203 11163 10232 11169
rect 10226 11160 10232 11163
rect 10284 11160 10290 11212
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 10796 11200 10824 11228
rect 10551 11172 10824 11200
rect 10965 11203 11023 11209
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 11072 11200 11100 11296
rect 12406 11268 12434 11296
rect 11440 11240 12434 11268
rect 11440 11209 11468 11240
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11072 11172 11253 11200
rect 10965 11163 11023 11169
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 9950 11132 9956 11144
rect 9784 11104 9956 11132
rect 9217 11095 9275 11101
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8570 11064 8576 11076
rect 8067 11036 8576 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 8665 11067 8723 11073
rect 8665 11033 8677 11067
rect 8711 11064 8723 11067
rect 9232 11064 9260 11095
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10980 11132 11008 11163
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11572 11172 11805 11200
rect 11572 11160 11578 11172
rect 11793 11169 11805 11172
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 10152 11104 11008 11132
rect 11057 11135 11115 11141
rect 8711 11036 9260 11064
rect 8711 11033 8723 11036
rect 8665 11027 8723 11033
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 10152 11064 10180 11104
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11698 11132 11704 11144
rect 11103 11104 11704 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12636 11132 12664 11308
rect 17402 11296 17408 11308
rect 17460 11296 17466 11348
rect 13354 11228 13360 11280
rect 13412 11228 13418 11280
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 14277 11271 14335 11277
rect 14277 11268 14289 11271
rect 13872 11240 14289 11268
rect 13872 11228 13878 11240
rect 14277 11237 14289 11240
rect 14323 11268 14335 11271
rect 15105 11271 15163 11277
rect 15105 11268 15117 11271
rect 14323 11240 15117 11268
rect 14323 11237 14335 11240
rect 14277 11231 14335 11237
rect 15105 11237 15117 11240
rect 15151 11268 15163 11271
rect 15286 11268 15292 11280
rect 15151 11240 15292 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 18141 11271 18199 11277
rect 18141 11237 18153 11271
rect 18187 11268 18199 11271
rect 18230 11268 18236 11280
rect 18187 11240 18236 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 18874 11228 18880 11280
rect 18932 11228 18938 11280
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 12802 11200 12808 11212
rect 12759 11172 12808 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 12986 11160 12992 11212
rect 13044 11160 13050 11212
rect 14001 11203 14059 11209
rect 14001 11200 14013 11203
rect 13188 11172 14013 11200
rect 12483 11104 12664 11132
rect 13004 11132 13032 11160
rect 13188 11132 13216 11172
rect 14001 11169 14013 11172
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14182 11160 14188 11212
rect 14240 11160 14246 11212
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 15194 11200 15200 11212
rect 14415 11172 15200 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 15194 11160 15200 11172
rect 15252 11200 15258 11212
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 15252 11172 15393 11200
rect 15252 11160 15258 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 16482 11160 16488 11212
rect 16540 11160 16546 11212
rect 17773 11203 17831 11209
rect 17773 11169 17785 11203
rect 17819 11169 17831 11203
rect 17773 11163 17831 11169
rect 13004 11104 13216 11132
rect 13265 11135 13323 11141
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 9640 11036 10180 11064
rect 9640 11024 9646 11036
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10594 11064 10600 11076
rect 10284 11036 10600 11064
rect 10284 11024 10290 11036
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 10686 11024 10692 11076
rect 10744 11024 10750 11076
rect 11606 11024 11612 11076
rect 11664 11064 11670 11076
rect 12529 11067 12587 11073
rect 12529 11064 12541 11067
rect 11664 11036 12541 11064
rect 11664 11024 11670 11036
rect 12529 11033 12541 11036
rect 12575 11033 12587 11067
rect 12529 11027 12587 11033
rect 12897 11067 12955 11073
rect 12897 11033 12909 11067
rect 12943 11064 12955 11067
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12943 11036 13093 11064
rect 12943 11033 12955 11036
rect 12897 11027 12955 11033
rect 13081 11033 13093 11036
rect 13127 11033 13139 11067
rect 13081 11027 13139 11033
rect 9858 10996 9864 11008
rect 7944 10968 9864 10996
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 10778 10996 10784 11008
rect 10192 10968 10784 10996
rect 10192 10956 10198 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 13280 10996 13308 11095
rect 13814 11024 13820 11076
rect 13872 11024 13878 11076
rect 13906 11024 13912 11076
rect 13964 11024 13970 11076
rect 14553 11067 14611 11073
rect 14553 11033 14565 11067
rect 14599 11064 14611 11067
rect 14826 11064 14832 11076
rect 14599 11036 14832 11064
rect 14599 11033 14611 11036
rect 14553 11027 14611 11033
rect 14826 11024 14832 11036
rect 14884 11064 14890 11076
rect 14936 11064 14964 11095
rect 15010 11092 15016 11144
rect 15068 11092 15074 11144
rect 17788 11073 17816 11163
rect 17773 11067 17831 11073
rect 14884 11036 15056 11064
rect 14884 11024 14890 11036
rect 13924 10996 13952 11024
rect 13280 10968 13952 10996
rect 14734 10956 14740 11008
rect 14792 10956 14798 11008
rect 15028 10996 15056 11036
rect 17773 11033 17785 11067
rect 17819 11064 17831 11067
rect 17862 11064 17868 11076
rect 17819 11036 17868 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 17126 10996 17132 11008
rect 15028 10968 17132 10996
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 1118 10752 1124 10804
rect 1176 10792 1182 10804
rect 1305 10795 1363 10801
rect 1305 10792 1317 10795
rect 1176 10764 1317 10792
rect 1176 10752 1182 10764
rect 1305 10761 1317 10764
rect 1351 10761 1363 10795
rect 1305 10755 1363 10761
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3200 10764 3249 10792
rect 3200 10752 3206 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 3237 10755 3295 10761
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 9306 10792 9312 10804
rect 6052 10764 9312 10792
rect 6052 10752 6058 10764
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 9456 10764 9628 10792
rect 9456 10752 9462 10764
rect 3326 10684 3332 10736
rect 3384 10684 3390 10736
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 8812 10696 9536 10724
rect 8812 10684 8818 10696
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 2464 10628 2789 10656
rect 2464 10616 2470 10628
rect 2777 10625 2789 10628
rect 2823 10625 2835 10659
rect 3510 10656 3516 10668
rect 2777 10619 2835 10625
rect 3252 10628 3516 10656
rect 1486 10548 1492 10600
rect 1544 10548 1550 10600
rect 1670 10548 1676 10600
rect 1728 10548 1734 10600
rect 3252 10597 3280 10628
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4212 10628 4261 10656
rect 4212 10616 4218 10628
rect 4249 10625 4261 10628
rect 4295 10656 4307 10659
rect 5810 10656 5816 10668
rect 4295 10628 5816 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 8386 10616 8392 10668
rect 8444 10616 8450 10668
rect 8588 10628 9444 10656
rect 8588 10600 8616 10628
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 1811 10560 2237 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 6546 10588 6552 10600
rect 5658 10560 6552 10588
rect 3237 10551 3295 10557
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 8570 10548 8576 10600
rect 8628 10548 8634 10600
rect 8662 10548 8668 10600
rect 8720 10548 8726 10600
rect 8846 10548 8852 10600
rect 8904 10548 8910 10600
rect 9416 10597 9444 10628
rect 9508 10597 9536 10696
rect 9600 10656 9628 10764
rect 10612 10764 10885 10792
rect 9784 10696 10088 10724
rect 9784 10656 9812 10696
rect 10060 10668 10088 10696
rect 10134 10684 10140 10736
rect 10192 10684 10198 10736
rect 9600 10628 9812 10656
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10557 9735 10591
rect 9784 10588 9812 10628
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 9916 10628 9996 10656
rect 9916 10616 9922 10628
rect 9968 10597 9996 10628
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 10152 10597 10180 10684
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10656 10379 10659
rect 10612 10656 10640 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11606 10792 11612 10804
rect 11011 10764 11612 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 11330 10724 11336 10736
rect 10827 10696 11336 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 13541 10727 13599 10733
rect 13541 10724 13553 10727
rect 12406 10696 13553 10724
rect 12406 10656 12434 10696
rect 13541 10693 13553 10696
rect 13587 10693 13599 10727
rect 13541 10687 13599 10693
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 13964 10696 14289 10724
rect 13964 10684 13970 10696
rect 14277 10693 14289 10696
rect 14323 10724 14335 10727
rect 14918 10724 14924 10736
rect 14323 10696 14924 10724
rect 14323 10693 14335 10696
rect 14277 10687 14335 10693
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 15488 10696 16344 10724
rect 10367 10628 10640 10656
rect 10796 10628 12434 10656
rect 13817 10659 13875 10665
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 10796 10600 10824 10628
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 15010 10656 15016 10668
rect 13863 10628 15016 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 15010 10616 15016 10628
rect 15068 10656 15074 10668
rect 15286 10656 15292 10668
rect 15068 10628 15292 10656
rect 15068 10616 15074 10628
rect 15286 10616 15292 10628
rect 15344 10656 15350 10668
rect 15488 10656 15516 10696
rect 15344 10628 15516 10656
rect 15344 10616 15350 10628
rect 9953 10591 10011 10597
rect 9784 10560 9878 10588
rect 9677 10551 9735 10557
rect 3513 10523 3571 10529
rect 3513 10489 3525 10523
rect 3559 10489 3571 10523
rect 3513 10483 3571 10489
rect 4525 10523 4583 10529
rect 4525 10489 4537 10523
rect 4571 10520 4583 10523
rect 4798 10520 4804 10532
rect 4571 10492 4804 10520
rect 4571 10489 4583 10492
rect 4525 10483 4583 10489
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 3528 10452 3556 10483
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 8680 10520 8708 10548
rect 9048 10520 9076 10551
rect 8680 10492 9076 10520
rect 3476 10424 3556 10452
rect 3476 10412 3482 10424
rect 8754 10412 8760 10464
rect 8812 10452 8818 10464
rect 8938 10452 8944 10464
rect 8812 10424 8944 10452
rect 8812 10412 8818 10424
rect 8938 10412 8944 10424
rect 8996 10452 9002 10464
rect 9692 10452 9720 10551
rect 9850 10529 9878 10560
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 9815 10523 9878 10529
rect 9815 10489 9827 10523
rect 9861 10492 9878 10523
rect 10045 10523 10103 10529
rect 9861 10489 9873 10492
rect 9815 10483 9873 10489
rect 10045 10489 10057 10523
rect 10091 10520 10103 10523
rect 10318 10520 10324 10532
rect 10091 10492 10324 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10520 10520 10548 10551
rect 10778 10548 10784 10600
rect 10836 10548 10842 10600
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 13998 10588 14004 10600
rect 13771 10560 14004 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 13832 10532 13860 10560
rect 13998 10548 14004 10560
rect 14056 10588 14062 10600
rect 14826 10588 14832 10600
rect 14056 10560 14832 10588
rect 14056 10548 14062 10560
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15194 10588 15200 10600
rect 14976 10560 15200 10588
rect 14976 10548 14982 10560
rect 15194 10548 15200 10560
rect 15252 10588 15258 10600
rect 15488 10597 15516 10628
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15620 10628 15853 10656
rect 15620 10616 15626 10628
rect 15841 10625 15853 10628
rect 15887 10656 15899 10659
rect 15887 10628 16160 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 16132 10597 16160 10628
rect 16316 10600 16344 10696
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10656 16451 10659
rect 16482 10656 16488 10668
rect 16439 10628 16488 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 17920 10628 18000 10656
rect 17920 10616 17926 10628
rect 17972 10600 18000 10628
rect 15473 10591 15531 10597
rect 15252 10560 15297 10588
rect 15252 10548 15258 10560
rect 15473 10557 15485 10591
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 16298 10548 16304 10600
rect 16356 10548 16362 10600
rect 17954 10548 17960 10600
rect 18012 10548 18018 10600
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10588 18291 10591
rect 18690 10588 18696 10600
rect 18279 10560 18696 10588
rect 18279 10557 18291 10560
rect 18233 10551 18291 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 18877 10591 18935 10597
rect 18877 10557 18889 10591
rect 18923 10588 18935 10591
rect 18923 10560 19104 10588
rect 18923 10557 18935 10560
rect 18877 10551 18935 10557
rect 10870 10520 10876 10532
rect 10520 10492 10876 10520
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 13814 10480 13820 10532
rect 13872 10480 13878 10532
rect 14182 10480 14188 10532
rect 14240 10520 14246 10532
rect 14277 10523 14335 10529
rect 14277 10520 14289 10523
rect 14240 10492 14289 10520
rect 14240 10480 14246 10492
rect 14277 10489 14289 10492
rect 14323 10489 14335 10523
rect 14277 10483 14335 10489
rect 8996 10424 9720 10452
rect 8996 10412 9002 10424
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10597 10455 10655 10461
rect 10597 10452 10609 10455
rect 10008 10424 10609 10452
rect 10008 10412 10014 10424
rect 10597 10421 10609 10424
rect 10643 10421 10655 10455
rect 10597 10415 10655 10421
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 14844 10452 14872 10548
rect 15565 10523 15623 10529
rect 15565 10489 15577 10523
rect 15611 10489 15623 10523
rect 15565 10483 15623 10489
rect 15102 10452 15108 10464
rect 14844 10424 15108 10452
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 15580 10452 15608 10483
rect 15930 10480 15936 10532
rect 15988 10480 15994 10532
rect 16206 10480 16212 10532
rect 16264 10520 16270 10532
rect 18325 10523 18383 10529
rect 18325 10520 18337 10523
rect 16264 10492 18337 10520
rect 16264 10480 16270 10492
rect 18325 10489 18337 10492
rect 18371 10489 18383 10523
rect 18325 10483 18383 10489
rect 19076 10464 19104 10560
rect 16482 10452 16488 10464
rect 15580 10424 16488 10452
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17460 10424 18061 10452
rect 17460 10412 17466 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18693 10455 18751 10461
rect 18693 10452 18705 10455
rect 18196 10424 18705 10452
rect 18196 10412 18202 10424
rect 18693 10421 18705 10424
rect 18739 10421 18751 10455
rect 18693 10415 18751 10421
rect 19058 10412 19064 10464
rect 19116 10412 19122 10464
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 3053 10251 3111 10257
rect 3053 10217 3065 10251
rect 3099 10248 3111 10251
rect 3142 10248 3148 10260
rect 3099 10220 3148 10248
rect 3099 10217 3111 10220
rect 3053 10211 3111 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 9950 10248 9956 10260
rect 9508 10220 9956 10248
rect 2590 10140 2596 10192
rect 2648 10180 2654 10192
rect 2777 10183 2835 10189
rect 2777 10180 2789 10183
rect 2648 10152 2789 10180
rect 2648 10140 2654 10152
rect 2777 10149 2789 10152
rect 2823 10149 2835 10183
rect 2777 10143 2835 10149
rect 3602 10140 3608 10192
rect 3660 10180 3666 10192
rect 7193 10183 7251 10189
rect 7193 10180 7205 10183
rect 3660 10152 7205 10180
rect 3660 10140 3666 10152
rect 7193 10149 7205 10152
rect 7239 10149 7251 10183
rect 7193 10143 7251 10149
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 9125 10183 9183 10189
rect 9125 10180 9137 10183
rect 7340 10152 9137 10180
rect 7340 10140 7346 10152
rect 9125 10149 9137 10152
rect 9171 10149 9183 10183
rect 9125 10143 9183 10149
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2961 10115 3019 10121
rect 2961 10112 2973 10115
rect 2556 10084 2973 10112
rect 2556 10072 2562 10084
rect 2961 10081 2973 10084
rect 3007 10081 3019 10115
rect 2961 10075 3019 10081
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 3234 10112 3240 10124
rect 3191 10084 3240 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 3375 10084 3525 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3513 10081 3525 10084
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 6641 10115 6699 10121
rect 6641 10081 6653 10115
rect 6687 10112 6699 10115
rect 8386 10112 8392 10124
rect 6687 10084 8392 10112
rect 6687 10081 6699 10084
rect 6641 10075 6699 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9048 10044 9076 10075
rect 9214 10072 9220 10124
rect 9272 10112 9278 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 9272 10084 9321 10112
rect 9272 10072 9278 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 9508 10044 9536 10220
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 11388 10220 12173 10248
rect 11388 10208 11394 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10217 12679 10251
rect 12621 10211 12679 10217
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 13814 10248 13820 10260
rect 12851 10220 13820 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 10652 10152 11008 10180
rect 10652 10140 10658 10152
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10112 10195 10115
rect 10226 10112 10232 10124
rect 10183 10084 10232 10112
rect 10183 10081 10195 10084
rect 10137 10075 10195 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 10318 10072 10324 10124
rect 10376 10072 10382 10124
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10870 10112 10876 10124
rect 10551 10084 10876 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 9048 10016 9536 10044
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 3510 9936 3516 9988
rect 3568 9976 3574 9988
rect 3697 9979 3755 9985
rect 3697 9976 3709 9979
rect 3568 9948 3709 9976
rect 3568 9936 3574 9948
rect 3697 9945 3709 9948
rect 3743 9976 3755 9979
rect 3878 9976 3884 9988
rect 3743 9948 3884 9976
rect 3743 9945 3755 9948
rect 3697 9939 3755 9945
rect 3878 9936 3884 9948
rect 3936 9936 3942 9988
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 6420 9880 6469 9908
rect 6420 9868 6426 9880
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6457 9871 6515 9877
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7926 9908 7932 9920
rect 7064 9880 7932 9908
rect 7064 9868 7070 9880
rect 7926 9868 7932 9880
rect 7984 9908 7990 9920
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 7984 9880 8493 9908
rect 7984 9868 7990 9880
rect 8481 9877 8493 9880
rect 8527 9877 8539 9911
rect 8481 9871 8539 9877
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 9585 9911 9643 9917
rect 9585 9908 9597 9911
rect 9539 9880 9597 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 9585 9877 9597 9880
rect 9631 9877 9643 9911
rect 9692 9908 9720 10007
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10428 10044 10456 10075
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10980 10121 11008 10152
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11238 10112 11244 10124
rect 11195 10084 11244 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 11572 10084 12357 10112
rect 11572 10072 11578 10084
rect 12345 10081 12357 10084
rect 12391 10112 12403 10115
rect 12434 10112 12440 10124
rect 12391 10084 12440 10112
rect 12391 10081 12403 10084
rect 12345 10075 12403 10081
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 12636 10112 12664 10211
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14240 10220 14289 10248
rect 14240 10208 14246 10220
rect 14277 10217 14289 10220
rect 14323 10248 14335 10251
rect 15194 10248 15200 10260
rect 14323 10220 15200 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15378 10208 15384 10260
rect 15436 10208 15442 10260
rect 15930 10208 15936 10260
rect 15988 10208 15994 10260
rect 15948 10180 15976 10208
rect 13096 10152 15976 10180
rect 12802 10112 12808 10124
rect 12636 10084 12808 10112
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 10100 10016 10456 10044
rect 12529 10047 12587 10053
rect 10100 10004 10106 10016
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 12618 10044 12624 10056
rect 12575 10016 12624 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 12618 10004 12624 10016
rect 12676 10044 12682 10056
rect 12986 10044 12992 10056
rect 12676 10016 12992 10044
rect 12676 10004 12682 10016
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10134 9976 10140 9988
rect 9999 9948 10140 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 10226 9936 10232 9988
rect 10284 9976 10290 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 10284 9948 10701 9976
rect 10284 9936 10290 9948
rect 10689 9945 10701 9948
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 10962 9908 10968 9920
rect 9692 9880 10968 9908
rect 9585 9871 9643 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11054 9868 11060 9920
rect 11112 9868 11118 9920
rect 11333 9911 11391 9917
rect 11333 9877 11345 9911
rect 11379 9908 11391 9911
rect 11698 9908 11704 9920
rect 11379 9880 11704 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12492 9880 12817 9908
rect 12492 9868 12498 9880
rect 12805 9877 12817 9880
rect 12851 9908 12863 9911
rect 13096 9908 13124 10152
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 13814 10112 13820 10124
rect 13771 10084 13820 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 14182 10072 14188 10124
rect 14240 10112 14246 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 14240 10084 14381 10112
rect 14240 10072 14246 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 15010 10072 15016 10124
rect 15068 10072 15074 10124
rect 15194 10072 15200 10124
rect 15252 10072 15258 10124
rect 14001 10047 14059 10053
rect 14001 10013 14013 10047
rect 14047 10013 14059 10047
rect 14001 10007 14059 10013
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 13449 9979 13507 9985
rect 13449 9976 13461 9979
rect 13219 9948 13461 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 13449 9945 13461 9948
rect 13495 9976 13507 9979
rect 13906 9976 13912 9988
rect 13495 9948 13912 9976
rect 13495 9945 13507 9948
rect 13449 9939 13507 9945
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 14016 9976 14044 10007
rect 14458 10004 14464 10056
rect 14516 10053 14522 10056
rect 14516 10047 14544 10053
rect 14532 10013 14544 10047
rect 15028 10044 15056 10072
rect 14516 10007 14544 10013
rect 14660 10016 15056 10044
rect 14516 10004 14522 10007
rect 14660 9976 14688 10016
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15396 10050 15516 10078
rect 15562 10072 15568 10124
rect 15620 10072 15626 10124
rect 15654 10072 15660 10124
rect 15712 10072 15718 10124
rect 15841 10115 15899 10121
rect 15841 10081 15853 10115
rect 15887 10112 15899 10115
rect 15948 10112 15976 10152
rect 16592 10152 17448 10180
rect 16592 10124 16620 10152
rect 15887 10084 15976 10112
rect 15887 10081 15899 10084
rect 15841 10075 15899 10081
rect 16482 10072 16488 10124
rect 16540 10072 16546 10124
rect 16574 10072 16580 10124
rect 16632 10072 16638 10124
rect 16758 10072 16764 10124
rect 16816 10072 16822 10124
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 17218 10112 17224 10124
rect 17175 10084 17224 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17420 10121 17448 10152
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10112 17463 10115
rect 17494 10112 17500 10124
rect 17451 10084 17500 10112
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18432 10084 18521 10112
rect 18432 10056 18460 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 15396 10044 15424 10050
rect 15160 10016 15424 10044
rect 15160 10004 15166 10016
rect 14016 9948 14688 9976
rect 15010 9936 15016 9988
rect 15068 9976 15074 9988
rect 15194 9976 15200 9988
rect 15068 9948 15200 9976
rect 15068 9936 15074 9948
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 12851 9880 13124 9908
rect 12851 9877 12863 9880
rect 12805 9871 12863 9877
rect 13262 9868 13268 9920
rect 13320 9868 13326 9920
rect 14642 9868 14648 9920
rect 14700 9868 14706 9920
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15105 9911 15163 9917
rect 15105 9908 15117 9911
rect 14976 9880 15117 9908
rect 14976 9868 14982 9880
rect 15105 9877 15117 9880
rect 15151 9877 15163 9911
rect 15488 9908 15516 10050
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 15580 10016 16313 10044
rect 15580 9988 15608 10016
rect 16301 10013 16313 10016
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 18414 10044 18420 10056
rect 18012 10016 18420 10044
rect 18012 10004 18018 10016
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 15562 9936 15568 9988
rect 15620 9936 15626 9988
rect 16114 9936 16120 9988
rect 16172 9976 16178 9988
rect 18506 9976 18512 9988
rect 16172 9948 18512 9976
rect 16172 9936 16178 9948
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 15488 9880 15761 9908
rect 15105 9871 15163 9877
rect 15749 9877 15761 9880
rect 15795 9877 15807 9911
rect 15749 9871 15807 9877
rect 15838 9868 15844 9920
rect 15896 9908 15902 9920
rect 16301 9911 16359 9917
rect 16301 9908 16313 9911
rect 15896 9880 16313 9908
rect 15896 9868 15902 9880
rect 16301 9877 16313 9880
rect 16347 9877 16359 9911
rect 16301 9871 16359 9877
rect 16390 9868 16396 9920
rect 16448 9868 16454 9920
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 18966 9908 18972 9920
rect 16899 9880 18972 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 8386 9664 8392 9716
rect 8444 9664 8450 9716
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10137 9707 10195 9713
rect 9916 9676 10088 9704
rect 9916 9664 9922 9676
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 1728 9608 3249 9636
rect 1728 9596 1734 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 10060 9636 10088 9676
rect 10137 9673 10149 9707
rect 10183 9704 10195 9707
rect 10594 9704 10600 9716
rect 10183 9676 10600 9704
rect 10183 9673 10195 9676
rect 10137 9667 10195 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 11020 9676 11529 9704
rect 11020 9664 11026 9676
rect 11517 9673 11529 9676
rect 11563 9673 11575 9707
rect 11517 9667 11575 9673
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9673 12495 9707
rect 12437 9667 12495 9673
rect 10060 9608 10640 9636
rect 3237 9599 3295 9605
rect 10612 9580 10640 9608
rect 10686 9596 10692 9648
rect 10744 9596 10750 9648
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 12345 9639 12403 9645
rect 10919 9608 12204 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5868 9540 6009 9568
rect 5868 9528 5874 9540
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6273 9571 6331 9577
rect 6273 9537 6285 9571
rect 6319 9568 6331 9571
rect 6362 9568 6368 9580
rect 6319 9540 6368 9568
rect 6319 9537 6331 9540
rect 6273 9531 6331 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 8754 9568 8760 9580
rect 7791 9540 8760 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 8754 9528 8760 9540
rect 8812 9568 8818 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8812 9540 8861 9568
rect 8812 9528 8818 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9122 9568 9128 9580
rect 9079 9540 9128 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2004 9472 2421 9500
rect 2004 9460 2010 9472
rect 2409 9469 2421 9472
rect 2455 9500 2467 9503
rect 2498 9500 2504 9512
rect 2455 9472 2504 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9500 2651 9503
rect 3142 9500 3148 9512
rect 2639 9472 3148 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 9048 9500 9076 9531
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9364 9540 9628 9568
rect 9364 9528 9370 9540
rect 8444 9472 9076 9500
rect 8444 9460 8450 9472
rect 9490 9460 9496 9512
rect 9548 9460 9554 9512
rect 9600 9509 9628 9540
rect 9784 9540 10548 9568
rect 9784 9509 9812 9540
rect 10520 9512 10548 9540
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10704 9568 10732 9596
rect 10704 9540 11008 9568
rect 9586 9503 9644 9509
rect 9586 9469 9598 9503
rect 9632 9469 9644 9503
rect 9586 9463 9644 9469
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 9999 9503 10057 9509
rect 9999 9469 10011 9503
rect 10045 9500 10057 9503
rect 10134 9500 10140 9512
rect 10045 9472 10140 9500
rect 10045 9469 10057 9472
rect 9999 9463 10057 9469
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10226 9460 10232 9512
rect 10284 9460 10290 9512
rect 10410 9509 10416 9512
rect 10377 9503 10416 9509
rect 10377 9469 10389 9503
rect 10377 9463 10416 9469
rect 10410 9460 10416 9463
rect 10468 9460 10474 9512
rect 10502 9460 10508 9512
rect 10560 9460 10566 9512
rect 10735 9503 10793 9509
rect 10735 9469 10747 9503
rect 10781 9500 10793 9503
rect 10870 9500 10876 9512
rect 10781 9472 10876 9500
rect 10781 9469 10793 9472
rect 10735 9463 10793 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 10980 9509 11008 9540
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11204 9540 11376 9568
rect 11204 9528 11210 9540
rect 11348 9512 11376 9540
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11480 9540 11836 9568
rect 11480 9528 11486 9540
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9469 11299 9503
rect 11241 9463 11299 9469
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 3421 9435 3479 9441
rect 3421 9432 3433 9435
rect 2823 9404 3433 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 3421 9401 3433 9404
rect 3467 9401 3479 9435
rect 3421 9395 3479 9401
rect 6730 9392 6736 9444
rect 6788 9392 6794 9444
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 9732 9404 9873 9432
rect 9732 9392 9738 9404
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 10597 9435 10655 9441
rect 10597 9432 10609 9435
rect 9861 9395 9919 9401
rect 10152 9404 10609 9432
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 3510 9364 3516 9376
rect 1636 9336 3516 9364
rect 1636 9324 1642 9336
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 7282 9364 7288 9376
rect 4304 9336 7288 9364
rect 4304 9324 4310 9336
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 8754 9324 8760 9376
rect 8812 9324 8818 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 10152 9364 10180 9404
rect 10597 9401 10609 9404
rect 10643 9401 10655 9435
rect 11256 9432 11284 9463
rect 11330 9460 11336 9512
rect 11388 9460 11394 9512
rect 11808 9509 11836 9540
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12176 9568 12204 9608
rect 12345 9605 12357 9639
rect 12391 9636 12403 9639
rect 12452 9636 12480 9667
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 14458 9704 14464 9716
rect 13044 9676 14464 9704
rect 13044 9664 13050 9676
rect 14458 9664 14464 9676
rect 14516 9704 14522 9716
rect 15654 9704 15660 9716
rect 14516 9676 15660 9704
rect 14516 9664 14522 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 18230 9664 18236 9716
rect 18288 9664 18294 9716
rect 18690 9664 18696 9716
rect 18748 9664 18754 9716
rect 12391 9608 12480 9636
rect 12391 9605 12403 9608
rect 12345 9599 12403 9605
rect 14090 9596 14096 9648
rect 14148 9636 14154 9648
rect 17681 9639 17739 9645
rect 17681 9636 17693 9639
rect 14148 9608 17693 9636
rect 14148 9596 14154 9608
rect 17681 9605 17693 9608
rect 17727 9605 17739 9639
rect 17681 9599 17739 9605
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18104 9608 18460 9636
rect 18104 9596 18110 9608
rect 11940 9540 12112 9568
rect 12176 9540 12480 9568
rect 11940 9528 11946 9540
rect 12084 9509 12112 9540
rect 12452 9509 12480 9540
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 12710 9568 12716 9580
rect 12636 9540 12716 9568
rect 11701 9503 11759 9509
rect 11701 9469 11713 9503
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 11794 9503 11852 9509
rect 11794 9469 11806 9503
rect 11840 9469 11852 9503
rect 11794 9463 11852 9469
rect 12069 9503 12127 9509
rect 12069 9469 12081 9503
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 12207 9503 12265 9509
rect 12207 9469 12219 9503
rect 12253 9500 12265 9503
rect 12437 9503 12495 9509
rect 12253 9472 12388 9500
rect 12253 9469 12265 9472
rect 12207 9463 12265 9469
rect 11606 9432 11612 9444
rect 11256 9404 11612 9432
rect 10597 9395 10655 9401
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 9180 9336 10180 9364
rect 11716 9364 11744 9463
rect 11977 9435 12035 9441
rect 11977 9401 11989 9435
rect 12023 9401 12035 9435
rect 12360 9432 12388 9472
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12636 9432 12664 9540
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 15194 9568 15200 9580
rect 12952 9540 14228 9568
rect 12952 9528 12958 9540
rect 12820 9432 12848 9528
rect 14200 9509 14228 9540
rect 14384 9540 15200 9568
rect 14384 9512 14412 9540
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15746 9528 15752 9580
rect 15804 9528 15810 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15948 9540 16037 9568
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14366 9460 14372 9512
rect 14424 9460 14430 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 12360 9404 12664 9432
rect 12728 9404 12848 9432
rect 11977 9395 12035 9401
rect 11790 9364 11796 9376
rect 11716 9336 11796 9364
rect 9180 9324 9186 9336
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 11992 9364 12020 9395
rect 12526 9364 12532 9376
rect 11992 9336 12532 9364
rect 12526 9324 12532 9336
rect 12584 9364 12590 9376
rect 12728 9364 12756 9404
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 14936 9432 14964 9463
rect 15102 9460 15108 9512
rect 15160 9509 15166 9512
rect 15160 9500 15172 9509
rect 15160 9472 15205 9500
rect 15160 9463 15172 9472
rect 15160 9460 15166 9463
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 15948 9509 15976 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 18138 9568 18144 9580
rect 16025 9531 16083 9537
rect 16408 9540 17632 9568
rect 16408 9512 16436 9540
rect 17604 9512 17632 9540
rect 17880 9540 18144 9568
rect 17880 9512 17908 9540
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15436 9472 15945 9500
rect 15436 9460 15442 9472
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 16390 9460 16396 9512
rect 16448 9460 16454 9512
rect 17497 9503 17555 9509
rect 17497 9469 17509 9503
rect 17543 9469 17555 9503
rect 17497 9463 17555 9469
rect 12952 9404 14964 9432
rect 17512 9432 17540 9463
rect 17586 9460 17592 9512
rect 17644 9460 17650 9512
rect 17678 9460 17684 9512
rect 17736 9460 17742 9512
rect 17862 9460 17868 9512
rect 17920 9460 17926 9512
rect 18432 9509 18460 9608
rect 18506 9528 18512 9580
rect 18564 9568 18570 9580
rect 19061 9571 19119 9577
rect 19061 9568 19073 9571
rect 18564 9540 19073 9568
rect 18564 9528 18570 9540
rect 19061 9537 19073 9540
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 17957 9503 18015 9509
rect 17957 9469 17969 9503
rect 18003 9469 18015 9503
rect 17957 9463 18015 9469
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 18417 9503 18475 9509
rect 18417 9469 18429 9503
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 17696 9432 17724 9460
rect 17512 9404 17724 9432
rect 12952 9392 12958 9404
rect 12584 9336 12756 9364
rect 12584 9324 12590 9336
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 17972 9364 18000 9463
rect 18248 9432 18276 9463
rect 18874 9460 18880 9512
rect 18932 9460 18938 9512
rect 18782 9432 18788 9444
rect 18248 9404 18788 9432
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 14976 9336 18000 9364
rect 14976 9324 14982 9336
rect 18138 9324 18144 9376
rect 18196 9324 18202 9376
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 2685 9163 2743 9169
rect 2685 9129 2697 9163
rect 2731 9160 2743 9163
rect 3142 9160 3148 9172
rect 2731 9132 3148 9160
rect 2731 9129 2743 9132
rect 2685 9123 2743 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 4246 9120 4252 9172
rect 4304 9120 4310 9172
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 4706 9160 4712 9172
rect 4387 9132 4712 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9160 4859 9163
rect 5537 9163 5595 9169
rect 4847 9132 5028 9160
rect 4847 9129 4859 9132
rect 4801 9123 4859 9129
rect 2406 9092 2412 9104
rect 2346 9064 2412 9092
rect 2406 9052 2412 9064
rect 2464 9052 2470 9104
rect 4264 9092 4292 9120
rect 2884 9064 4292 9092
rect 4525 9095 4583 9101
rect 2884 9033 2912 9064
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 4724 9092 4752 9120
rect 4571 9064 4660 9092
rect 4724 9064 4936 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 4632 9036 4660 9064
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2746 8996 2881 9024
rect 842 8916 848 8968
rect 900 8916 906 8968
rect 1118 8916 1124 8968
rect 1176 8916 1182 8968
rect 2746 8956 2774 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 3789 9027 3847 9033
rect 3789 8993 3801 9027
rect 3835 9024 3847 9027
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3835 8996 4077 9024
rect 3835 8993 3847 8996
rect 3789 8987 3847 8993
rect 4065 8993 4077 8996
rect 4111 9024 4123 9027
rect 4154 9024 4160 9036
rect 4111 8996 4160 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4614 8984 4620 9036
rect 4672 8984 4678 9036
rect 4908 9033 4936 9064
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 2608 8928 2774 8956
rect 3053 8959 3111 8965
rect 2608 8832 2636 8928
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 2590 8780 2596 8832
rect 2648 8780 2654 8832
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 3068 8820 3096 8919
rect 3510 8916 3516 8968
rect 3568 8956 3574 8968
rect 4706 8956 4712 8968
rect 3568 8928 4712 8956
rect 3568 8916 3574 8928
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 3697 8891 3755 8897
rect 3697 8857 3709 8891
rect 3743 8888 3755 8891
rect 4617 8891 4675 8897
rect 4617 8888 4629 8891
rect 3743 8860 4629 8888
rect 3743 8857 3755 8860
rect 3697 8851 3755 8857
rect 4617 8857 4629 8860
rect 4663 8857 4675 8891
rect 5000 8888 5028 9132
rect 5537 9129 5549 9163
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 5552 9092 5580 9123
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 6236 9132 7573 9160
rect 6236 9120 6242 9132
rect 7561 9129 7573 9132
rect 7607 9160 7619 9163
rect 8665 9163 8723 9169
rect 7607 9132 8340 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 6089 9095 6147 9101
rect 6089 9092 6101 9095
rect 5552 9064 6101 9092
rect 6089 9061 6101 9064
rect 6135 9061 6147 9095
rect 6089 9055 6147 9061
rect 6730 9052 6736 9104
rect 6788 9052 6794 9104
rect 8312 9101 8340 9132
rect 8665 9129 8677 9163
rect 8711 9160 8723 9163
rect 8846 9160 8852 9172
rect 8711 9132 8852 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 9548 9132 10333 9160
rect 9548 9120 9554 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 11330 9120 11336 9172
rect 11388 9120 11394 9172
rect 11440 9132 11744 9160
rect 8297 9095 8355 9101
rect 8297 9061 8309 9095
rect 8343 9092 8355 9095
rect 9582 9092 9588 9104
rect 8343 9064 9588 9092
rect 8343 9061 8355 9064
rect 8297 9055 8355 9061
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 9953 9095 10011 9101
rect 9953 9061 9965 9095
rect 9999 9092 10011 9095
rect 10410 9092 10416 9104
rect 9999 9064 10416 9092
rect 9999 9061 10011 9064
rect 9953 9055 10011 9061
rect 10410 9052 10416 9064
rect 10468 9052 10474 9104
rect 10870 9052 10876 9104
rect 10928 9092 10934 9104
rect 11440 9101 11468 9132
rect 10965 9095 11023 9101
rect 10965 9092 10977 9095
rect 10928 9064 10977 9092
rect 10928 9052 10934 9064
rect 10965 9061 10977 9064
rect 11011 9061 11023 9095
rect 10965 9055 11023 9061
rect 11165 9095 11223 9101
rect 11165 9061 11177 9095
rect 11211 9092 11223 9095
rect 11425 9095 11483 9101
rect 11211 9064 11376 9092
rect 11211 9061 11223 9064
rect 11165 9055 11223 9061
rect 5350 8984 5356 9036
rect 5408 8984 5414 9036
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 8812 8996 9689 9024
rect 8812 8984 8818 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 9835 9027 9893 9033
rect 9835 8993 9847 9027
rect 9881 9024 9893 9027
rect 10045 9027 10103 9033
rect 9881 8993 9904 9024
rect 9835 8987 9904 8993
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 9024 10195 9027
rect 10318 9024 10324 9036
rect 10183 8996 10324 9024
rect 10183 8993 10195 8996
rect 10137 8987 10195 8993
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 4617 8851 4675 8857
rect 4724 8860 5028 8888
rect 8036 8888 8064 8919
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8168 8928 8217 8956
rect 8168 8916 8174 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8294 8888 8300 8900
rect 8036 8860 8300 8888
rect 2740 8792 3096 8820
rect 2740 8780 2746 8792
rect 3602 8780 3608 8832
rect 3660 8780 3666 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 3936 8792 4353 8820
rect 3936 8780 3942 8792
rect 4341 8789 4353 8792
rect 4387 8820 4399 8823
rect 4724 8820 4752 8860
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 4387 8792 4752 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 9766 8820 9772 8832
rect 4856 8792 9772 8820
rect 4856 8780 4862 8792
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9876 8820 9904 8987
rect 10060 8888 10088 8987
rect 10318 8984 10324 8996
rect 10376 9024 10382 9036
rect 11180 9024 11208 9055
rect 10376 8996 11208 9024
rect 11348 9024 11376 9064
rect 11425 9061 11437 9095
rect 11471 9061 11483 9095
rect 11425 9055 11483 9061
rect 11514 9052 11520 9104
rect 11572 9092 11578 9104
rect 11625 9095 11683 9101
rect 11625 9092 11637 9095
rect 11572 9064 11637 9092
rect 11572 9052 11578 9064
rect 11625 9061 11637 9064
rect 11671 9061 11683 9095
rect 11716 9092 11744 9132
rect 11790 9120 11796 9172
rect 11848 9120 11854 9172
rect 12802 9120 12808 9172
rect 12860 9120 12866 9172
rect 14458 9120 14464 9172
rect 14516 9160 14522 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 14516 9132 15761 9160
rect 14516 9120 14522 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 12158 9092 12164 9104
rect 11716 9064 12164 9092
rect 11625 9055 11683 9061
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 12820 9092 12848 9120
rect 12820 9064 14964 9092
rect 11532 9024 11560 9052
rect 11348 8996 11560 9024
rect 10376 8984 10382 8996
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 14090 9024 14096 9036
rect 13412 8996 14096 9024
rect 13412 8984 13418 8996
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 14274 8984 14280 9036
rect 14332 8984 14338 9036
rect 14936 9033 14964 9064
rect 15562 9052 15568 9104
rect 15620 9052 15626 9104
rect 16301 9095 16359 9101
rect 16301 9061 16313 9095
rect 16347 9092 16359 9095
rect 16390 9092 16396 9104
rect 16347 9064 16396 9092
rect 16347 9061 16359 9064
rect 16301 9055 16359 9061
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 14369 9027 14427 9033
rect 14369 8993 14381 9027
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 12710 8956 12716 8968
rect 10928 8928 12716 8956
rect 10928 8916 10934 8928
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 12768 8928 13553 8956
rect 12768 8916 12774 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 14001 8959 14059 8965
rect 14001 8925 14013 8959
rect 14047 8956 14059 8959
rect 14384 8956 14412 8987
rect 14458 8956 14464 8968
rect 14047 8928 14464 8956
rect 14047 8925 14059 8928
rect 14001 8919 14059 8925
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 10060 8860 11192 8888
rect 10778 8820 10784 8832
rect 9876 8792 10784 8820
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11164 8829 11192 8860
rect 11790 8848 11796 8900
rect 11848 8888 11854 8900
rect 12158 8888 12164 8900
rect 11848 8860 12164 8888
rect 11848 8848 11854 8860
rect 12158 8848 12164 8860
rect 12216 8888 12222 8900
rect 13817 8891 13875 8897
rect 13817 8888 13829 8891
rect 12216 8860 13829 8888
rect 12216 8848 12222 8860
rect 13817 8857 13829 8860
rect 13863 8857 13875 8891
rect 14568 8888 14596 8987
rect 15010 8984 15016 9036
rect 15068 8984 15074 9036
rect 15102 8984 15108 9036
rect 15160 8984 15166 9036
rect 15654 8984 15660 9036
rect 15712 8984 15718 9036
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 8993 15899 9027
rect 15841 8987 15899 8993
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 9024 16635 9027
rect 16758 9024 16764 9036
rect 16623 8996 16764 9024
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 14829 8959 14887 8965
rect 14829 8925 14841 8959
rect 14875 8956 14887 8959
rect 15028 8956 15056 8984
rect 14875 8928 15056 8956
rect 14875 8925 14887 8928
rect 14829 8919 14887 8925
rect 15120 8888 15148 8984
rect 14568 8860 15148 8888
rect 15856 8888 15884 8987
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 17218 9024 17224 9036
rect 17083 8996 17224 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 17862 9024 17868 9036
rect 17451 8996 17868 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 18414 8916 18420 8968
rect 18472 8956 18478 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 18472 8928 18521 8956
rect 18472 8916 18478 8928
rect 18509 8925 18521 8928
rect 18555 8956 18567 8959
rect 18616 8956 18644 8987
rect 18555 8928 18644 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 16482 8888 16488 8900
rect 15856 8860 16488 8888
rect 13817 8851 13875 8857
rect 16482 8848 16488 8860
rect 16540 8888 16546 8900
rect 18598 8888 18604 8900
rect 16540 8860 18604 8888
rect 16540 8848 16546 8860
rect 18598 8848 18604 8860
rect 18656 8848 18662 8900
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11195 8792 11621 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 11609 8789 11621 8792
rect 11655 8820 11667 8823
rect 13262 8820 13268 8832
rect 11655 8792 13268 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 16114 8820 16120 8832
rect 14231 8792 16120 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 1118 8576 1124 8628
rect 1176 8616 1182 8628
rect 1489 8619 1547 8625
rect 1489 8616 1501 8619
rect 1176 8588 1501 8616
rect 1176 8576 1182 8588
rect 1489 8585 1501 8588
rect 1535 8585 1547 8619
rect 1489 8579 1547 8585
rect 3500 8619 3558 8625
rect 3500 8585 3512 8619
rect 3546 8616 3558 8619
rect 3602 8616 3608 8628
rect 3546 8588 3608 8616
rect 3546 8585 3558 8588
rect 3500 8579 3558 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5408 8588 5733 8616
rect 5408 8576 5414 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8251 8588 8984 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 1581 8551 1639 8557
rect 1581 8517 1593 8551
rect 1627 8548 1639 8551
rect 2041 8551 2099 8557
rect 2041 8548 2053 8551
rect 1627 8520 2053 8548
rect 1627 8517 1639 8520
rect 1581 8511 1639 8517
rect 2041 8517 2053 8520
rect 2087 8517 2099 8551
rect 2041 8511 2099 8517
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 4985 8551 5043 8557
rect 4985 8548 4997 8551
rect 4672 8520 4997 8548
rect 4672 8508 4678 8520
rect 4985 8517 4997 8520
rect 5031 8548 5043 8551
rect 8754 8548 8760 8560
rect 5031 8520 8760 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 8956 8548 8984 8588
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9088 8588 9505 8616
rect 9088 8576 9094 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 11146 8576 11152 8628
rect 11204 8576 11210 8628
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 12066 8576 12072 8628
rect 12124 8576 12130 8628
rect 18322 8616 18328 8628
rect 13188 8588 18328 8616
rect 11164 8548 11192 8576
rect 8956 8520 11192 8548
rect 842 8440 848 8492
rect 900 8480 906 8492
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 900 8452 3249 8480
rect 900 8440 906 8452
rect 3237 8449 3249 8452
rect 3283 8480 3295 8483
rect 3283 8452 5856 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 5828 8424 5856 8452
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 6822 8480 6828 8492
rect 6411 8452 6828 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 8294 8480 8300 8492
rect 7699 8452 8300 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8294 8440 8300 8452
rect 8352 8480 8358 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8352 8452 8861 8480
rect 8352 8440 8358 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11992 8480 12020 8576
rect 12161 8483 12219 8489
rect 12161 8480 12173 8483
rect 11112 8452 11652 8480
rect 11992 8452 12173 8480
rect 11112 8440 11118 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1578 8412 1584 8424
rect 1443 8384 1584 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 1765 8375 1823 8381
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8412 2099 8415
rect 2590 8412 2596 8424
rect 2087 8384 2596 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 1780 8276 1808 8375
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 5810 8372 5816 8424
rect 5868 8372 5874 8424
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8412 6147 8415
rect 7282 8412 7288 8424
rect 6135 8384 7288 8412
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7834 8372 7840 8424
rect 7892 8372 7898 8424
rect 9122 8372 9128 8424
rect 9180 8372 9186 8424
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 10376 8384 11437 8412
rect 10376 8372 10382 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 11514 8372 11520 8424
rect 11572 8372 11578 8424
rect 11624 8412 11652 8452
rect 12161 8449 12173 8452
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12452 8452 12848 8480
rect 12452 8424 12480 8452
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11624 8384 11713 8412
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 2498 8344 2504 8356
rect 1912 8316 2504 8344
rect 1912 8304 1918 8316
rect 2498 8304 2504 8316
rect 2556 8304 2562 8356
rect 2746 8316 4002 8344
rect 1946 8276 1952 8288
rect 1780 8248 1952 8276
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 2746 8276 2774 8316
rect 6914 8304 6920 8356
rect 6972 8304 6978 8356
rect 7745 8347 7803 8353
rect 7745 8313 7757 8347
rect 7791 8344 7803 8347
rect 8018 8344 8024 8356
rect 7791 8316 8024 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 10870 8344 10876 8356
rect 8220 8316 10876 8344
rect 2464 8248 2774 8276
rect 6932 8276 6960 8304
rect 8220 8276 8248 8316
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11146 8344 11152 8356
rect 11020 8316 11152 8344
rect 11020 8304 11026 8316
rect 11146 8304 11152 8316
rect 11204 8344 11210 8356
rect 11808 8344 11836 8375
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 11940 8384 12357 8412
rect 11940 8372 11946 8384
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12434 8372 12440 8424
rect 12492 8372 12498 8424
rect 12820 8421 12848 8452
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8381 12679 8415
rect 12621 8375 12679 8381
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 11204 8316 11836 8344
rect 11977 8347 12035 8353
rect 11204 8304 11210 8316
rect 11977 8313 11989 8347
rect 12023 8344 12035 8347
rect 12069 8347 12127 8353
rect 12069 8344 12081 8347
rect 12023 8316 12081 8344
rect 12023 8313 12035 8316
rect 11977 8307 12035 8313
rect 12069 8313 12081 8316
rect 12115 8313 12127 8347
rect 12069 8307 12127 8313
rect 12158 8304 12164 8356
rect 12216 8344 12222 8356
rect 12636 8344 12664 8375
rect 12986 8372 12992 8424
rect 13044 8372 13050 8424
rect 13188 8421 13216 8588
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 13357 8551 13415 8557
rect 13357 8517 13369 8551
rect 13403 8548 13415 8551
rect 16574 8548 16580 8560
rect 13403 8520 16580 8548
rect 13403 8517 13415 8520
rect 13357 8511 13415 8517
rect 16574 8508 16580 8520
rect 16632 8548 16638 8560
rect 18414 8548 18420 8560
rect 16632 8520 16988 8548
rect 16632 8508 16638 8520
rect 13998 8480 14004 8492
rect 13740 8452 14004 8480
rect 13740 8421 13768 8452
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8480 14887 8483
rect 14875 8452 15148 8480
rect 14875 8449 14887 8452
rect 14829 8443 14887 8449
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 12216 8316 12664 8344
rect 13004 8344 13032 8372
rect 13740 8344 13768 8375
rect 13906 8372 13912 8424
rect 13964 8372 13970 8424
rect 14185 8415 14243 8421
rect 14185 8381 14197 8415
rect 14231 8412 14243 8415
rect 14274 8412 14280 8424
rect 14231 8384 14280 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 13004 8316 13768 8344
rect 12216 8304 12222 8316
rect 6932 8248 8248 8276
rect 2464 8236 2470 8248
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9033 8279 9091 8285
rect 9033 8276 9045 8279
rect 8812 8248 9045 8276
rect 8812 8236 8818 8248
rect 9033 8245 9045 8248
rect 9079 8245 9091 8279
rect 9033 8239 9091 8245
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 12434 8276 12440 8288
rect 11480 8248 12440 8276
rect 11480 8236 11486 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 12526 8236 12532 8288
rect 12584 8236 12590 8288
rect 12897 8279 12955 8285
rect 12897 8245 12909 8279
rect 12943 8276 12955 8279
rect 12986 8276 12992 8288
rect 12943 8248 12992 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 14200 8276 14228 8375
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14752 8344 14780 8440
rect 14415 8316 14780 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14844 8276 14872 8443
rect 15120 8424 15148 8452
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 16960 8489 16988 8520
rect 17926 8520 18420 8548
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17770 8440 17776 8492
rect 17828 8480 17834 8492
rect 17926 8480 17954 8520
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 18874 8508 18880 8560
rect 18932 8548 18938 8560
rect 18932 8520 19104 8548
rect 18932 8508 18938 8520
rect 19076 8489 19104 8520
rect 17828 8452 17954 8480
rect 19061 8483 19119 8489
rect 17828 8440 17834 8452
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 15102 8372 15108 8424
rect 15160 8372 15166 8424
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 15749 8415 15807 8421
rect 15252 8384 15277 8412
rect 15252 8372 15258 8384
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 16206 8412 16212 8424
rect 15795 8384 16212 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16390 8372 16396 8424
rect 16448 8372 16454 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 17420 8412 17448 8440
rect 16899 8384 17448 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17644 8384 18061 8412
rect 17644 8372 17650 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 18877 8415 18935 8421
rect 18877 8381 18889 8415
rect 18923 8381 18935 8415
rect 18877 8375 18935 8381
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 15212 8344 15240 8372
rect 16408 8344 16436 8372
rect 15068 8316 16436 8344
rect 15068 8304 15074 8316
rect 17862 8304 17868 8356
rect 17920 8344 17926 8356
rect 18892 8344 18920 8375
rect 17920 8316 18920 8344
rect 17920 8304 17926 8316
rect 14200 8248 14872 8276
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 18230 8276 18236 8288
rect 15344 8248 18236 8276
rect 15344 8236 15350 8248
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 18690 8236 18696 8288
rect 18748 8236 18754 8288
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 1854 8032 1860 8084
rect 1912 8032 1918 8084
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 7006 8072 7012 8084
rect 2004 8044 7012 8072
rect 2004 8032 2010 8044
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7432 8044 7573 8072
rect 7432 8032 7438 8044
rect 7561 8041 7573 8044
rect 7607 8072 7619 8075
rect 7834 8072 7840 8084
rect 7607 8044 7840 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 8389 8075 8447 8081
rect 8036 8044 8340 8072
rect 1578 7964 1584 8016
rect 1636 8004 1642 8016
rect 1673 8007 1731 8013
rect 1673 8004 1685 8007
rect 1636 7976 1685 8004
rect 1636 7964 1642 7976
rect 1673 7973 1685 7976
rect 1719 7973 1731 8007
rect 1673 7967 1731 7973
rect 1964 7945 1992 8032
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7905 2007 7939
rect 1949 7899 2007 7905
rect 5442 7896 5448 7948
rect 5500 7896 5506 7948
rect 5810 7896 5816 7948
rect 5868 7896 5874 7948
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 8036 7945 8064 8044
rect 8110 7964 8116 8016
rect 8168 7964 8174 8016
rect 8312 8004 8340 8044
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8478 8072 8484 8084
rect 8435 8044 8484 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 9033 8075 9091 8081
rect 8680 8044 8892 8072
rect 8570 8004 8576 8016
rect 8312 7976 8576 8004
rect 8570 7964 8576 7976
rect 8628 8004 8634 8016
rect 8680 8013 8708 8044
rect 8665 8007 8723 8013
rect 8665 8004 8677 8007
rect 8628 7976 8677 8004
rect 8628 7964 8634 7976
rect 8665 7973 8677 7976
rect 8711 7973 8723 8007
rect 8665 7967 8723 7973
rect 8754 7964 8760 8016
rect 8812 7964 8818 8016
rect 8864 8004 8892 8044
rect 9033 8041 9045 8075
rect 9079 8072 9091 8075
rect 10226 8072 10232 8084
rect 9079 8044 10232 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 11992 8044 16344 8072
rect 10778 8004 10784 8016
rect 8864 7976 10784 8004
rect 10778 7964 10784 7976
rect 10836 7964 10842 8016
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 11992 8004 12020 8044
rect 11572 7976 12020 8004
rect 12268 7976 16252 8004
rect 11572 7964 11578 7976
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7300 7908 7849 7936
rect 7300 7880 7328 7908
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7905 8079 7939
rect 8229 7939 8287 7945
rect 8229 7936 8241 7939
rect 8021 7899 8079 7905
rect 8220 7905 8241 7936
rect 8275 7905 8287 7939
rect 8220 7899 8287 7905
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5644 7840 6101 7868
rect 5644 7809 5672 7840
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 8220 7868 8248 7899
rect 8478 7896 8484 7948
rect 8536 7896 8542 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9398 7936 9404 7948
rect 8904 7908 9404 7936
rect 8904 7896 8910 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10502 7936 10508 7948
rect 9824 7908 10508 7936
rect 9824 7896 9830 7908
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11698 7936 11704 7948
rect 11296 7908 11704 7936
rect 11296 7896 11302 7908
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11809 7945 11837 7976
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 12158 7896 12164 7948
rect 12216 7896 12222 7948
rect 12268 7945 12296 7976
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 12434 7896 12440 7948
rect 12492 7896 12498 7948
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7936 12679 7939
rect 12986 7936 12992 7948
rect 12667 7908 12992 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 13170 7896 13176 7948
rect 13228 7896 13234 7948
rect 13630 7896 13636 7948
rect 13688 7896 13694 7948
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 13780 7908 14197 7936
rect 13780 7896 13786 7908
rect 14185 7905 14197 7908
rect 14231 7936 14243 7939
rect 15010 7936 15016 7948
rect 14231 7908 15016 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7905 15439 7939
rect 15381 7899 15439 7905
rect 8864 7868 8892 7896
rect 8220 7840 8892 7868
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10410 7868 10416 7880
rect 10284 7840 10416 7868
rect 10284 7828 10290 7840
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 12452 7868 12480 7896
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12452 7840 12725 7868
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 5629 7803 5687 7809
rect 5629 7769 5641 7803
rect 5675 7769 5687 7803
rect 12434 7800 12440 7812
rect 5629 7763 5687 7769
rect 7116 7772 12440 7800
rect 1670 7692 1676 7744
rect 1728 7692 1734 7744
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 7116 7732 7144 7772
rect 12434 7760 12440 7772
rect 12492 7760 12498 7812
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 12820 7800 12848 7831
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 13004 7868 13032 7896
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13004 7840 14289 7868
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 15396 7868 15424 7899
rect 15930 7896 15936 7948
rect 15988 7896 15994 7948
rect 14277 7831 14335 7837
rect 14384 7840 15424 7868
rect 14384 7812 14412 7840
rect 13630 7800 13636 7812
rect 12676 7772 13636 7800
rect 12676 7760 12682 7772
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 13998 7760 14004 7812
rect 14056 7800 14062 7812
rect 14366 7800 14372 7812
rect 14056 7772 14372 7800
rect 14056 7760 14062 7772
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 14550 7760 14556 7812
rect 14608 7760 14614 7812
rect 15010 7760 15016 7812
rect 15068 7760 15074 7812
rect 16224 7800 16252 7976
rect 16316 7945 16344 8044
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18598 8072 18604 8084
rect 18472 8044 18604 8072
rect 18472 8032 18478 8044
rect 18598 8032 18604 8044
rect 18656 8072 18662 8084
rect 18656 8044 18828 8072
rect 18656 8032 18662 8044
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 16390 7896 16396 7948
rect 16448 7896 16454 7948
rect 16574 7896 16580 7948
rect 16632 7896 16638 7948
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17644 7908 17693 7936
rect 17644 7896 17650 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 18230 7896 18236 7948
rect 18288 7896 18294 7948
rect 18506 7896 18512 7948
rect 18564 7896 18570 7948
rect 18800 7945 18828 8044
rect 18785 7939 18843 7945
rect 18785 7905 18797 7939
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 18966 7896 18972 7948
rect 19024 7896 19030 7948
rect 18601 7871 18659 7877
rect 18601 7868 18613 7871
rect 16684 7840 18613 7868
rect 16684 7800 16712 7840
rect 18601 7837 18613 7840
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 16224 7772 16712 7800
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 17828 7772 17877 7800
rect 17828 7760 17834 7772
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 4120 7704 7144 7732
rect 4120 7692 4126 7704
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 10410 7732 10416 7744
rect 9732 7704 10416 7732
rect 9732 7692 9738 7704
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 11238 7692 11244 7744
rect 11296 7692 11302 7744
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 13078 7732 13084 7744
rect 12032 7704 13084 7732
rect 12032 7692 12038 7704
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 16117 7735 16175 7741
rect 16117 7732 16129 7735
rect 13504 7704 16129 7732
rect 13504 7692 13510 7704
rect 16117 7701 16129 7704
rect 16163 7701 16175 7735
rect 16117 7695 16175 7701
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2556 7500 2605 7528
rect 2556 7488 2562 7500
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 2593 7491 2651 7497
rect 842 7352 848 7404
rect 900 7352 906 7404
rect 2406 7324 2412 7336
rect 2254 7296 2412 7324
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 1118 7216 1124 7268
rect 1176 7216 1182 7268
rect 2608 7256 2636 7491
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 5868 7500 6193 7528
rect 5868 7488 5874 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 6181 7491 6239 7497
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 10318 7528 10324 7540
rect 8987 7500 10324 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 11698 7488 11704 7540
rect 11756 7488 11762 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 11931 7500 13400 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 5460 7460 5488 7488
rect 6733 7463 6791 7469
rect 6733 7460 6745 7463
rect 5460 7432 6745 7460
rect 6733 7429 6745 7432
rect 6779 7429 6791 7463
rect 6733 7423 6791 7429
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 7064 7432 9996 7460
rect 7064 7420 7070 7432
rect 4154 7352 4160 7404
rect 4212 7352 4218 7404
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6880 7364 7297 7392
rect 6880 7352 6886 7364
rect 7285 7361 7297 7364
rect 7331 7392 7343 7395
rect 8846 7392 8852 7404
rect 7331 7364 7972 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 4172 7324 4200 7352
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 4172 7296 4261 7324
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 4249 7287 4307 7293
rect 4816 7296 7113 7324
rect 2958 7256 2964 7268
rect 2608 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7256 3022 7268
rect 4816 7256 4844 7296
rect 7101 7293 7113 7296
rect 7147 7324 7159 7327
rect 7147 7296 7696 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 3016 7228 4844 7256
rect 4893 7259 4951 7265
rect 3016 7216 3022 7228
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 7558 7256 7564 7268
rect 4939 7228 7564 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 3786 7148 3792 7200
rect 3844 7148 3850 7200
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 4246 7188 4252 7200
rect 4203 7160 4252 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 4246 7148 4252 7160
rect 4304 7188 4310 7200
rect 6914 7188 6920 7200
rect 4304 7160 6920 7188
rect 4304 7148 4310 7160
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7193 7191 7251 7197
rect 7193 7157 7205 7191
rect 7239 7188 7251 7191
rect 7374 7188 7380 7200
rect 7239 7160 7380 7188
rect 7239 7157 7251 7160
rect 7193 7151 7251 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7668 7188 7696 7296
rect 7944 7256 7972 7364
rect 8036 7364 8708 7392
rect 8036 7336 8064 7364
rect 8018 7284 8024 7336
rect 8076 7284 8082 7336
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8168 7296 8401 7324
rect 8168 7284 8174 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 8680 7333 8708 7364
rect 8772 7364 8852 7392
rect 8772 7333 8800 7364
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9732 7364 9873 7392
rect 9732 7352 9738 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9968 7392 9996 7432
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9968 7364 10333 7392
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 9766 7324 9772 7336
rect 8757 7287 8815 7293
rect 9692 7296 9772 7324
rect 9306 7256 9312 7268
rect 7944 7228 9312 7256
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 9692 7265 9720 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 9968 7333 9996 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 11716 7392 11744 7488
rect 13372 7472 13400 7500
rect 13556 7500 14047 7528
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 12584 7432 13124 7460
rect 12584 7420 12590 7432
rect 11716 7364 11928 7392
rect 10321 7355 10379 7361
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10137 7327 10195 7333
rect 10137 7293 10149 7327
rect 10183 7324 10195 7327
rect 10226 7324 10232 7336
rect 10183 7296 10232 7324
rect 10183 7293 10195 7296
rect 10137 7287 10195 7293
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 11330 7324 11336 7336
rect 10827 7296 11336 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 11422 7284 11428 7336
rect 11480 7284 11486 7336
rect 11698 7284 11704 7336
rect 11756 7284 11762 7336
rect 11790 7284 11796 7336
rect 11848 7284 11854 7336
rect 11900 7324 11928 7364
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 11900 7296 12449 7324
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7293 12679 7327
rect 12621 7287 12679 7293
rect 13096 7320 13124 7432
rect 13354 7420 13360 7472
rect 13412 7420 13418 7472
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13556 7392 13584 7500
rect 13722 7420 13728 7472
rect 13780 7420 13786 7472
rect 13311 7364 13584 7392
rect 14019 7392 14047 7500
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 18690 7528 18696 7540
rect 14148 7500 18696 7528
rect 14148 7488 14154 7500
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 18874 7488 18880 7540
rect 18932 7488 18938 7540
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 18046 7460 18052 7472
rect 14608 7432 18052 7460
rect 14608 7420 14614 7432
rect 14019 7364 15056 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13173 7327 13231 7333
rect 13173 7320 13185 7327
rect 13096 7293 13185 7320
rect 13219 7293 13231 7327
rect 13096 7292 13231 7293
rect 13173 7287 13231 7292
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7326 13599 7327
rect 13587 7324 13743 7326
rect 14090 7324 14096 7336
rect 13587 7298 14096 7324
rect 13587 7293 13599 7298
rect 13715 7296 14096 7298
rect 13541 7287 13599 7293
rect 9677 7259 9735 7265
rect 9677 7225 9689 7259
rect 9723 7225 9735 7259
rect 10873 7259 10931 7265
rect 9677 7219 9735 7225
rect 9876 7228 10824 7256
rect 9876 7188 9904 7228
rect 7668 7160 9904 7188
rect 9953 7191 10011 7197
rect 9953 7157 9965 7191
rect 9999 7188 10011 7191
rect 10226 7188 10232 7200
rect 9999 7160 10232 7188
rect 9999 7157 10011 7160
rect 9953 7151 10011 7157
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10468 7160 10701 7188
rect 10468 7148 10474 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10796 7188 10824 7228
rect 10873 7225 10885 7259
rect 10919 7256 10931 7259
rect 11146 7256 11152 7268
rect 10919 7228 11152 7256
rect 10919 7225 10931 7228
rect 10873 7219 10931 7225
rect 11146 7216 11152 7228
rect 11204 7256 11210 7268
rect 11808 7256 11836 7284
rect 11204 7228 11836 7256
rect 11204 7216 11210 7228
rect 12066 7216 12072 7268
rect 12124 7216 12130 7268
rect 11054 7188 11060 7200
rect 10796 7160 11060 7188
rect 10689 7151 10747 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11514 7148 11520 7200
rect 11572 7148 11578 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12636 7188 12664 7287
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 14274 7284 14280 7336
rect 14332 7284 14338 7336
rect 13262 7216 13268 7268
rect 13320 7256 13326 7268
rect 13817 7259 13875 7265
rect 13817 7256 13829 7259
rect 13320 7228 13829 7256
rect 13320 7216 13326 7228
rect 13817 7225 13829 7228
rect 13863 7225 13875 7259
rect 15028 7256 15056 7364
rect 15120 7333 15148 7432
rect 18046 7420 18052 7432
rect 18104 7420 18110 7472
rect 18138 7420 18144 7472
rect 18196 7420 18202 7472
rect 18322 7420 18328 7472
rect 18380 7420 18386 7472
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 17770 7392 17776 7404
rect 15436 7364 17776 7392
rect 15436 7352 15442 7364
rect 17770 7352 17776 7364
rect 17828 7392 17834 7404
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17828 7364 17969 7392
rect 17828 7352 17834 7364
rect 17957 7361 17969 7364
rect 18003 7392 18015 7395
rect 18003 7364 18092 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7324 15807 7327
rect 15838 7324 15844 7336
rect 15795 7296 15844 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 16080 7296 16865 7324
rect 16080 7284 16086 7296
rect 16853 7293 16865 7296
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 17678 7324 17684 7336
rect 16991 7296 17684 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 18064 7333 18092 7364
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18156 7324 18184 7420
rect 18340 7392 18368 7420
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 18340 7364 18705 7392
rect 18693 7361 18705 7364
rect 18739 7361 18751 7395
rect 18892 7392 18920 7488
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18892 7364 19073 7392
rect 18693 7355 18751 7361
rect 18874 7324 18880 7336
rect 18156 7296 18880 7324
rect 18049 7287 18107 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 18230 7256 18236 7268
rect 15028 7228 18236 7256
rect 13817 7219 13875 7225
rect 18230 7216 18236 7228
rect 18288 7216 18294 7268
rect 11756 7160 12664 7188
rect 11756 7148 11762 7160
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 18690 7188 18696 7200
rect 13136 7160 18696 7188
rect 13136 7148 13142 7160
rect 18690 7148 18696 7160
rect 18748 7188 18754 7200
rect 18984 7188 19012 7364
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 18748 7160 19012 7188
rect 18748 7148 18754 7160
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 1946 6944 1952 6996
rect 2004 6944 2010 6996
rect 4062 6984 4068 6996
rect 3804 6956 4068 6984
rect 1670 6808 1676 6860
rect 1728 6808 1734 6860
rect 1857 6851 1915 6857
rect 1857 6817 1869 6851
rect 1903 6848 1915 6851
rect 1964 6848 1992 6944
rect 3804 6925 3832 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 4154 6944 4160 6996
rect 4212 6944 4218 6996
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 10229 6987 10287 6993
rect 7248 6956 7420 6984
rect 7248 6944 7254 6956
rect 3589 6919 3647 6925
rect 3589 6885 3601 6919
rect 3635 6916 3647 6919
rect 3789 6919 3847 6925
rect 3635 6885 3648 6916
rect 3589 6879 3648 6885
rect 3789 6885 3801 6919
rect 3835 6885 3847 6919
rect 4172 6916 4200 6944
rect 5258 6916 5264 6928
rect 3789 6879 3847 6885
rect 3988 6888 5264 6916
rect 1903 6820 1992 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 2958 6808 2964 6860
rect 3016 6808 3022 6860
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3283 6820 3464 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 1118 6740 1124 6792
rect 1176 6780 1182 6792
rect 1489 6783 1547 6789
rect 1489 6780 1501 6783
rect 1176 6752 1501 6780
rect 1176 6740 1182 6752
rect 1489 6749 1501 6752
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 1995 6752 2329 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2317 6749 2329 6752
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 3436 6721 3464 6820
rect 3620 6780 3648 6879
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 3988 6848 4016 6888
rect 5258 6876 5264 6888
rect 5316 6876 5322 6928
rect 3927 6820 4016 6848
rect 4065 6851 4123 6857
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4338 6848 4344 6860
rect 4111 6820 4344 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4338 6808 4344 6820
rect 4396 6848 4402 6860
rect 5350 6848 5356 6860
rect 4396 6820 5356 6848
rect 4396 6808 4402 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 7392 6834 7420 6956
rect 10229 6953 10241 6987
rect 10275 6984 10287 6987
rect 10410 6984 10416 6996
rect 10275 6956 10416 6984
rect 10275 6953 10287 6956
rect 10229 6947 10287 6953
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 10560 6956 11468 6984
rect 10560 6944 10566 6956
rect 10042 6876 10048 6928
rect 10100 6916 10106 6928
rect 11440 6916 11468 6956
rect 11606 6944 11612 6996
rect 11664 6944 11670 6996
rect 15562 6984 15568 6996
rect 13372 6956 15568 6984
rect 11790 6916 11796 6928
rect 10100 6888 10732 6916
rect 10100 6876 10106 6888
rect 7926 6808 7932 6860
rect 7984 6808 7990 6860
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6817 10379 6851
rect 10704 6848 10732 6888
rect 11440 6888 11796 6916
rect 11330 6848 11336 6860
rect 10704 6820 11336 6848
rect 10321 6811 10379 6817
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3620 6752 3985 6780
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 3421 6715 3479 6721
rect 3421 6681 3433 6715
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 4982 6712 4988 6724
rect 4856 6684 4988 6712
rect 4856 6672 4862 6684
rect 4982 6672 4988 6684
rect 5040 6672 5046 6724
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 3053 6647 3111 6653
rect 3053 6644 3065 6647
rect 2556 6616 3065 6644
rect 2556 6604 2562 6616
rect 3053 6613 3065 6616
rect 3099 6613 3111 6647
rect 3053 6607 3111 6613
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3786 6644 3792 6656
rect 3651 6616 3792 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5442 6644 5448 6656
rect 4948 6616 5448 6644
rect 4948 6604 4954 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6012 6644 6040 6743
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8294 6780 8300 6792
rect 7791 6752 8300 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8294 6740 8300 6752
rect 8352 6780 8358 6792
rect 8754 6780 8760 6792
rect 8352 6752 8760 6780
rect 8352 6740 8358 6752
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 10336 6780 10364 6811
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 10336 6752 10916 6780
rect 9692 6712 9720 6740
rect 10045 6715 10103 6721
rect 10045 6712 10057 6715
rect 9692 6684 10057 6712
rect 10045 6681 10057 6684
rect 10091 6681 10103 6715
rect 10045 6675 10103 6681
rect 10888 6656 10916 6752
rect 11146 6740 11152 6792
rect 11204 6740 11210 6792
rect 7374 6644 7380 6656
rect 6012 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6644 7438 6656
rect 9398 6644 9404 6656
rect 7432 6616 9404 6644
rect 7432 6604 7438 6616
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 10870 6604 10876 6656
rect 10928 6604 10934 6656
rect 11164 6644 11192 6740
rect 11440 6721 11468 6888
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 12268 6888 12480 6916
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 11664 6820 11713 6848
rect 11664 6808 11670 6820
rect 11701 6817 11713 6820
rect 11747 6817 11759 6851
rect 11701 6811 11759 6817
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6848 11943 6851
rect 12268 6848 12296 6888
rect 11931 6820 12296 6848
rect 11931 6817 11943 6820
rect 11885 6811 11943 6817
rect 12342 6808 12348 6860
rect 12400 6808 12406 6860
rect 12452 6848 12480 6888
rect 12526 6848 12532 6860
rect 12452 6820 12532 6848
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 12952 6820 13277 6848
rect 12952 6808 12958 6820
rect 13265 6817 13277 6820
rect 13311 6848 13323 6851
rect 13372 6848 13400 6956
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 13814 6916 13820 6928
rect 13311 6820 13400 6848
rect 13715 6888 13820 6916
rect 13311 6817 13323 6820
rect 13265 6811 13323 6817
rect 13715 6789 13743 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15194 6916 15200 6928
rect 14424 6888 15200 6916
rect 14424 6876 14430 6888
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 16758 6916 16764 6928
rect 15396 6888 16764 6916
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 15286 6848 15292 6860
rect 14231 6820 15292 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 13700 6783 13758 6789
rect 11900 6752 13584 6780
rect 11900 6724 11928 6752
rect 11425 6715 11483 6721
rect 11425 6681 11437 6715
rect 11471 6681 11483 6715
rect 11425 6675 11483 6681
rect 11882 6672 11888 6724
rect 11940 6672 11946 6724
rect 12161 6715 12219 6721
rect 12161 6681 12173 6715
rect 12207 6712 12219 6715
rect 12802 6712 12808 6724
rect 12207 6684 12808 6712
rect 12207 6681 12219 6684
rect 12161 6675 12219 6681
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 13446 6712 13452 6724
rect 12912 6684 13452 6712
rect 11606 6644 11612 6656
rect 11164 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11756 6616 11805 6644
rect 11756 6604 11762 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12912 6644 12940 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 13556 6721 13584 6752
rect 13700 6749 13712 6783
rect 13746 6749 13758 6783
rect 13700 6743 13758 6749
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 13998 6780 14004 6792
rect 13955 6752 14004 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6681 13599 6715
rect 13541 6675 13599 6681
rect 12400 6616 12940 6644
rect 12400 6604 12406 6616
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13832 6644 13860 6743
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 13228 6616 13860 6644
rect 14384 6644 14412 6743
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 15396 6780 15424 6888
rect 15838 6808 15844 6860
rect 15896 6808 15902 6860
rect 16408 6857 16436 6888
rect 16758 6876 16764 6888
rect 16816 6916 16822 6928
rect 17586 6916 17592 6928
rect 16816 6888 17592 6916
rect 16816 6876 16822 6888
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 16393 6851 16451 6857
rect 16393 6817 16405 6851
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 16850 6808 16856 6860
rect 16908 6808 16914 6860
rect 17221 6851 17279 6857
rect 17221 6817 17233 6851
rect 17267 6848 17279 6851
rect 18138 6848 18144 6860
rect 17267 6820 18144 6848
rect 17267 6817 17279 6820
rect 17221 6811 17279 6817
rect 15160 6752 15424 6780
rect 15160 6740 15166 6752
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 17236 6780 17264 6811
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 18598 6808 18604 6860
rect 18656 6808 18662 6860
rect 15528 6752 17264 6780
rect 17497 6783 17555 6789
rect 15528 6740 15534 6752
rect 17497 6749 17509 6783
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 15378 6672 15384 6724
rect 15436 6712 15442 6724
rect 15657 6715 15715 6721
rect 15657 6712 15669 6715
rect 15436 6684 15669 6712
rect 15436 6672 15442 6684
rect 15657 6681 15669 6684
rect 15703 6712 15715 6715
rect 15746 6712 15752 6724
rect 15703 6684 15752 6712
rect 15703 6681 15715 6684
rect 15657 6675 15715 6681
rect 15746 6672 15752 6684
rect 15804 6672 15810 6724
rect 16022 6712 16028 6724
rect 15856 6684 16028 6712
rect 15856 6644 15884 6684
rect 16022 6672 16028 6684
rect 16080 6672 16086 6724
rect 16390 6672 16396 6724
rect 16448 6672 16454 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 17512 6712 17540 6743
rect 17770 6740 17776 6792
rect 17828 6740 17834 6792
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 17926 6752 18521 6780
rect 16816 6684 17540 6712
rect 17788 6712 17816 6740
rect 17926 6712 17954 6752
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 17788 6684 17954 6712
rect 16816 6672 16822 6684
rect 14384 6616 15884 6644
rect 13228 6604 13234 6616
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16574 6644 16580 6656
rect 15988 6616 16580 6644
rect 15988 6604 15994 6616
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 17218 6644 17224 6656
rect 16908 6616 17224 6644
rect 16908 6604 16914 6616
rect 17218 6604 17224 6616
rect 17276 6644 17282 6656
rect 17954 6644 17960 6656
rect 17276 6616 17960 6644
rect 17276 6604 17282 6616
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 4028 6412 4261 6440
rect 4028 6400 4034 6412
rect 4249 6409 4261 6412
rect 4295 6440 4307 6443
rect 4338 6440 4344 6452
rect 4295 6412 4344 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 4982 6400 4988 6452
rect 5040 6400 5046 6452
rect 6086 6400 6092 6452
rect 6144 6400 6150 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6328 6412 6469 6440
rect 6328 6400 6334 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 6457 6403 6515 6409
rect 6564 6412 11621 6440
rect 4847 6375 4905 6381
rect 4847 6341 4859 6375
rect 4893 6372 4905 6375
rect 4893 6344 5672 6372
rect 4893 6341 4905 6344
rect 4847 6335 4905 6341
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 5644 6313 5672 6344
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 5316 6276 5365 6304
rect 5316 6264 5322 6276
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 6104 6304 6132 6400
rect 5675 6276 6132 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4264 6208 4537 6236
rect 3970 6128 3976 6180
rect 4028 6128 4034 6180
rect 4062 6128 4068 6180
rect 4120 6128 4126 6180
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 4264 6177 4292 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 4985 6233 5043 6239
rect 4985 6199 4997 6233
rect 5031 6230 5043 6233
rect 5074 6230 5080 6248
rect 5031 6202 5080 6230
rect 5031 6199 5043 6202
rect 4985 6193 5043 6199
rect 5074 6196 5080 6202
rect 5132 6196 5138 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 5276 6208 5457 6236
rect 4264 6171 4323 6177
rect 4264 6168 4277 6171
rect 4212 6140 4277 6168
rect 4212 6128 4218 6140
rect 4265 6137 4277 6140
rect 4311 6137 4323 6171
rect 4265 6131 4323 6137
rect 4356 6140 4752 6168
rect 3988 6100 4016 6128
rect 4356 6100 4384 6140
rect 3988 6072 4384 6100
rect 4430 6060 4436 6112
rect 4488 6060 4494 6112
rect 4614 6060 4620 6112
rect 4672 6060 4678 6112
rect 4724 6109 4752 6140
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6069 4767 6103
rect 5276 6100 5304 6208
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6564 6236 6592 6412
rect 11609 6409 11621 6412
rect 11655 6409 11667 6443
rect 11609 6403 11667 6409
rect 13633 6443 13691 6449
rect 13633 6409 13645 6443
rect 13679 6440 13691 6443
rect 13814 6440 13820 6452
rect 13679 6412 13820 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 14182 6400 14188 6452
rect 14240 6400 14246 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 17494 6440 17500 6452
rect 15712 6412 17500 6440
rect 15712 6400 15718 6412
rect 17494 6400 17500 6412
rect 17552 6440 17558 6452
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 17552 6412 17693 6440
rect 17552 6400 17558 6412
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 17681 6403 17739 6409
rect 18230 6400 18236 6452
rect 18288 6400 18294 6452
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6341 6883 6375
rect 8757 6375 8815 6381
rect 6825 6335 6883 6341
rect 7484 6344 8432 6372
rect 6227 6208 6592 6236
rect 6641 6239 6699 6245
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 6840 6236 6868 6335
rect 7484 6313 7512 6344
rect 8404 6316 8432 6344
rect 8757 6341 8769 6375
rect 8803 6341 8815 6375
rect 8757 6335 8815 6341
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8386 6264 8392 6316
rect 8444 6264 8450 6316
rect 6687 6208 6868 6236
rect 7285 6239 7343 6245
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 8312 6236 8340 6264
rect 7331 6208 8340 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 5350 6128 5356 6180
rect 5408 6168 5414 6180
rect 5552 6168 5580 6199
rect 8478 6196 8484 6248
rect 8536 6196 8542 6248
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6236 8631 6239
rect 8772 6236 8800 6335
rect 11330 6332 11336 6384
rect 11388 6372 11394 6384
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 11388 6344 11529 6372
rect 11388 6332 11394 6344
rect 11517 6341 11529 6344
rect 11563 6341 11575 6375
rect 11517 6335 11575 6341
rect 12618 6332 12624 6384
rect 12676 6332 12682 6384
rect 18598 6372 18604 6384
rect 15166 6344 16804 6372
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 9180 6276 9229 6304
rect 9180 6264 9186 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9456 6276 9781 6304
rect 9456 6264 9462 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6304 10103 6307
rect 10134 6304 10140 6316
rect 10091 6276 10140 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13265 6307 13323 6313
rect 13265 6304 13277 6307
rect 13228 6276 13277 6304
rect 13228 6264 13234 6276
rect 13265 6273 13277 6276
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 15166 6304 15194 6344
rect 16776 6316 16804 6344
rect 16868 6344 18604 6372
rect 14332 6276 15194 6304
rect 14332 6264 14338 6276
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16022 6304 16028 6316
rect 15979 6276 16028 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16758 6264 16764 6316
rect 16816 6264 16822 6316
rect 8619 6208 8800 6236
rect 11793 6239 11851 6245
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6236 12035 6239
rect 12023 6208 12388 6236
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 7193 6171 7251 6177
rect 7193 6168 7205 6171
rect 5408 6140 7205 6168
rect 5408 6128 5414 6140
rect 7193 6137 7205 6140
rect 7239 6168 7251 6171
rect 8496 6168 8524 6196
rect 7239 6140 8524 6168
rect 9125 6171 9183 6177
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 9125 6137 9137 6171
rect 9171 6168 9183 6171
rect 10042 6168 10048 6180
rect 9171 6140 10048 6168
rect 9171 6137 9183 6140
rect 9125 6131 9183 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10502 6168 10508 6180
rect 10152 6140 10508 6168
rect 5442 6100 5448 6112
rect 5276 6072 5448 6100
rect 4709 6063 4767 6069
rect 5442 6060 5448 6072
rect 5500 6100 5506 6112
rect 6454 6100 6460 6112
rect 5500 6072 6460 6100
rect 5500 6060 5506 6072
rect 6454 6060 6460 6072
rect 6512 6060 6518 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 8352 6072 8401 6100
rect 8352 6060 8358 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 9490 6100 9496 6112
rect 8628 6072 9496 6100
rect 8628 6060 8634 6072
rect 9490 6060 9496 6072
rect 9548 6100 9554 6112
rect 10152 6100 10180 6140
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 11808 6168 11836 6199
rect 12253 6171 12311 6177
rect 12253 6168 12265 6171
rect 11808 6140 12265 6168
rect 9548 6072 10180 6100
rect 9548 6060 9554 6072
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 11808 6100 11836 6140
rect 12253 6137 12265 6140
rect 12299 6137 12311 6171
rect 12360 6168 12388 6208
rect 12894 6196 12900 6248
rect 12952 6196 12958 6248
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 12437 6171 12495 6177
rect 12437 6168 12449 6171
rect 12360 6140 12449 6168
rect 12253 6131 12311 6137
rect 12437 6137 12449 6140
rect 12483 6168 12495 6171
rect 12526 6168 12532 6180
rect 12483 6140 12532 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 10928 6072 11836 6100
rect 12268 6100 12296 6131
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12802 6128 12808 6180
rect 12860 6128 12866 6180
rect 12912 6100 12940 6196
rect 13004 6112 13032 6199
rect 12268 6072 12940 6100
rect 10928 6060 10934 6072
rect 12986 6060 12992 6112
rect 13044 6060 13050 6112
rect 13096 6100 13124 6199
rect 13354 6196 13360 6248
rect 13412 6196 13418 6248
rect 13538 6196 13544 6248
rect 13596 6196 13602 6248
rect 14060 6239 14118 6245
rect 14060 6205 14072 6239
rect 14106 6236 14118 6239
rect 14366 6236 14372 6248
rect 14106 6208 14372 6236
rect 14106 6205 14118 6208
rect 13832 6180 13978 6202
rect 14060 6199 14118 6205
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 14458 6196 14464 6248
rect 14516 6196 14522 6248
rect 15838 6236 15844 6248
rect 15166 6208 15844 6236
rect 13814 6128 13820 6180
rect 13872 6177 13978 6180
rect 13872 6174 13994 6177
rect 13872 6128 13878 6174
rect 13936 6171 13994 6174
rect 13936 6137 13948 6171
rect 13982 6137 13994 6171
rect 14476 6168 14504 6196
rect 15166 6168 15194 6208
rect 15838 6196 15844 6208
rect 15896 6236 15902 6248
rect 16868 6236 16896 6344
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 15896 6208 16896 6236
rect 15896 6196 15902 6208
rect 16960 6180 16988 6267
rect 17052 6245 17080 6344
rect 18598 6332 18604 6344
rect 18656 6332 18662 6384
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 18322 6304 18328 6316
rect 17552 6276 18328 6304
rect 17552 6264 17558 6276
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 18690 6264 18696 6316
rect 18748 6264 18754 6316
rect 17037 6239 17095 6245
rect 17037 6205 17049 6239
rect 17083 6205 17095 6239
rect 17770 6236 17776 6248
rect 17037 6199 17095 6205
rect 17144 6208 17776 6236
rect 14476 6140 15194 6168
rect 13936 6131 13994 6137
rect 15746 6128 15752 6180
rect 15804 6168 15810 6180
rect 16942 6168 16948 6180
rect 15804 6140 16948 6168
rect 15804 6128 15810 6140
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 17144 6100 17172 6208
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 17954 6196 17960 6248
rect 18012 6196 18018 6248
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 17586 6128 17592 6180
rect 17644 6128 17650 6180
rect 13096 6072 17172 6100
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 18248 6100 18276 6199
rect 18414 6196 18420 6248
rect 18472 6196 18478 6248
rect 18782 6196 18788 6248
rect 18840 6236 18846 6248
rect 18877 6239 18935 6245
rect 18877 6236 18889 6239
rect 18840 6208 18889 6236
rect 18840 6196 18846 6208
rect 18877 6205 18889 6208
rect 18923 6205 18935 6239
rect 18877 6199 18935 6205
rect 17276 6072 18276 6100
rect 17276 6060 17282 6072
rect 18414 6060 18420 6112
rect 18472 6100 18478 6112
rect 18800 6100 18828 6196
rect 18472 6072 18828 6100
rect 18472 6060 18478 6072
rect 19058 6060 19064 6112
rect 19116 6060 19122 6112
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 2464 5868 3648 5896
rect 2464 5856 2470 5868
rect 2498 5788 2504 5840
rect 2556 5788 2562 5840
rect 842 5720 848 5772
rect 900 5760 906 5772
rect 2225 5763 2283 5769
rect 2225 5760 2237 5763
rect 900 5732 2237 5760
rect 900 5720 906 5732
rect 2225 5729 2237 5732
rect 2271 5729 2283 5763
rect 2225 5723 2283 5729
rect 3620 5624 3648 5868
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 4430 5856 4436 5908
rect 4488 5856 4494 5908
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 4856 5868 5396 5896
rect 4856 5856 4862 5868
rect 4356 5769 4384 5856
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4448 5760 4476 5856
rect 4816 5800 5304 5828
rect 4816 5769 4844 5800
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4448 5732 4629 5760
rect 4341 5723 4399 5729
rect 4617 5729 4629 5732
rect 4663 5729 4675 5763
rect 4617 5723 4675 5729
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 4632 5692 4660 5723
rect 5276 5701 5304 5800
rect 5368 5769 5396 5868
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 8570 5896 8576 5908
rect 6788 5868 7880 5896
rect 6788 5856 6794 5868
rect 7852 5828 7880 5868
rect 8312 5868 8576 5896
rect 8312 5828 8340 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 9272 5868 9413 5896
rect 9272 5856 9278 5868
rect 9401 5865 9413 5868
rect 9447 5865 9459 5899
rect 9401 5859 9459 5865
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 10870 5896 10876 5908
rect 10459 5868 10876 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11514 5896 11520 5908
rect 11072 5868 11520 5896
rect 7852 5800 8418 5828
rect 9582 5788 9588 5840
rect 9640 5828 9646 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 9640 5800 10977 5828
rect 9640 5788 9646 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 10965 5791 11023 5797
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 6641 5763 6699 5769
rect 6641 5760 6653 5763
rect 5592 5732 6653 5760
rect 5592 5720 5598 5732
rect 6641 5729 6653 5732
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 7282 5720 7288 5772
rect 7340 5720 7346 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7432 5732 7665 5760
rect 7432 5720 7438 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10321 5763 10379 5769
rect 9723 5732 9996 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 4632 5664 5089 5692
rect 5077 5661 5089 5664
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5307 5664 5825 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 4798 5624 4804 5636
rect 3620 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 5184 5624 5212 5655
rect 6454 5652 6460 5704
rect 6512 5692 6518 5704
rect 6914 5692 6920 5704
rect 6512 5664 6920 5692
rect 6512 5652 6518 5664
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 5040 5596 7205 5624
rect 5040 5584 5046 5596
rect 7193 5593 7205 5596
rect 7239 5593 7251 5627
rect 7193 5587 7251 5593
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 4893 5559 4951 5565
rect 4893 5556 4905 5559
rect 4488 5528 4905 5556
rect 4488 5516 4494 5528
rect 4893 5525 4905 5528
rect 4939 5525 4951 5559
rect 7300 5556 7328 5720
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8294 5692 8300 5704
rect 7975 5664 8300 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 9968 5633 9996 5732
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 11072 5760 11100 5868
rect 11514 5856 11520 5868
rect 11572 5896 11578 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 11572 5868 12633 5896
rect 11572 5856 11578 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 15470 5896 15476 5908
rect 12621 5859 12679 5865
rect 13648 5868 15476 5896
rect 11149 5831 11207 5837
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 11422 5828 11428 5840
rect 11195 5800 11428 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 13648 5828 13676 5868
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15620 5868 15669 5896
rect 15620 5856 15626 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 17678 5856 17684 5908
rect 17736 5896 17742 5908
rect 18969 5899 19027 5905
rect 18969 5896 18981 5899
rect 17736 5868 18981 5896
rect 17736 5856 17742 5868
rect 18969 5865 18981 5868
rect 19015 5865 19027 5899
rect 18969 5859 19027 5865
rect 11532 5800 12204 5828
rect 11532 5769 11560 5800
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 10367 5732 11345 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5760 11667 5763
rect 11974 5760 11980 5772
rect 11655 5732 11980 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 10410 5652 10416 5704
rect 10468 5692 10474 5704
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 10468 5664 10517 5692
rect 10468 5652 10474 5664
rect 10505 5661 10517 5664
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11624 5692 11652 5723
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 11020 5664 11652 5692
rect 11020 5652 11026 5664
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11848 5664 12081 5692
rect 11848 5652 11854 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 9585 5627 9643 5633
rect 9585 5624 9597 5627
rect 9364 5596 9597 5624
rect 9364 5584 9370 5596
rect 9585 5593 9597 5596
rect 9631 5593 9643 5627
rect 9585 5587 9643 5593
rect 9953 5627 10011 5633
rect 9953 5593 9965 5627
rect 9999 5593 10011 5627
rect 12176 5624 12204 5800
rect 13556 5800 13676 5828
rect 15764 5800 15976 5828
rect 12342 5720 12348 5772
rect 12400 5720 12406 5772
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5760 12495 5763
rect 12710 5760 12716 5772
rect 12483 5732 12716 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 13556 5769 13584 5800
rect 13449 5763 13507 5769
rect 13449 5729 13461 5763
rect 13495 5729 13507 5763
rect 13449 5723 13507 5729
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 13354 5692 13360 5704
rect 12851 5664 13360 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 13464 5692 13492 5723
rect 13630 5720 13636 5772
rect 13688 5720 13694 5772
rect 13817 5763 13875 5769
rect 13817 5729 13829 5763
rect 13863 5760 13875 5763
rect 14090 5760 14096 5772
rect 13863 5732 14096 5760
rect 13863 5729 13875 5732
rect 13817 5723 13875 5729
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5760 14427 5763
rect 15378 5760 15384 5772
rect 14415 5732 15384 5760
rect 14415 5729 14427 5732
rect 14369 5723 14427 5729
rect 13648 5692 13676 5720
rect 13464 5664 13676 5692
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 14384 5692 14412 5723
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 15764 5769 15792 5800
rect 15948 5772 15976 5800
rect 18598 5788 18604 5840
rect 18656 5788 18662 5840
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 15838 5720 15844 5772
rect 15896 5720 15902 5772
rect 15930 5720 15936 5772
rect 15988 5720 15994 5772
rect 16390 5720 16396 5772
rect 16448 5760 16454 5772
rect 17218 5760 17224 5772
rect 16448 5732 17224 5760
rect 16448 5720 16454 5732
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18506 5760 18512 5772
rect 18003 5732 18512 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 13771 5664 14412 5692
rect 14461 5695 14519 5701
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14461 5661 14473 5695
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15519 5664 16129 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 13265 5627 13323 5633
rect 13265 5624 13277 5627
rect 12176 5596 13277 5624
rect 9953 5587 10011 5593
rect 13265 5593 13277 5596
rect 13311 5624 13323 5627
rect 14476 5624 14504 5655
rect 15746 5624 15752 5636
rect 13311 5596 13952 5624
rect 14476 5596 15752 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 7926 5556 7932 5568
rect 7300 5528 7932 5556
rect 4893 5519 4951 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 11793 5559 11851 5565
rect 11793 5525 11805 5559
rect 11839 5556 11851 5559
rect 12710 5556 12716 5568
rect 11839 5528 12716 5556
rect 11839 5525 11851 5528
rect 11793 5519 11851 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13722 5556 13728 5568
rect 13044 5528 13728 5556
rect 13044 5516 13050 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 13924 5556 13952 5596
rect 15746 5584 15752 5596
rect 15804 5584 15810 5636
rect 15194 5556 15200 5568
rect 13924 5528 15200 5556
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15856 5556 15884 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 17972 5692 18000 5723
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 18874 5720 18880 5772
rect 18932 5720 18938 5772
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 16356 5664 18000 5692
rect 16356 5652 16362 5664
rect 18046 5652 18052 5704
rect 18104 5692 18110 5704
rect 18966 5692 18972 5704
rect 18104 5664 18972 5692
rect 18104 5652 18110 5664
rect 18966 5652 18972 5664
rect 19024 5692 19030 5704
rect 19076 5692 19104 5723
rect 19024 5664 19104 5692
rect 19024 5652 19030 5664
rect 16942 5584 16948 5636
rect 17000 5624 17006 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 17000 5596 17417 5624
rect 17000 5584 17006 5596
rect 17405 5593 17417 5596
rect 17451 5624 17463 5627
rect 18506 5624 18512 5636
rect 17451 5596 18512 5624
rect 17451 5593 17463 5596
rect 17405 5587 17463 5593
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 16114 5556 16120 5568
rect 15344 5528 16120 5556
rect 15344 5516 15350 5528
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 3684 5355 3742 5361
rect 3684 5321 3696 5355
rect 3730 5352 3742 5355
rect 4154 5352 4160 5364
rect 3730 5324 4160 5352
rect 3730 5321 3742 5324
rect 3684 5315 3742 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 5000 5324 5457 5352
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 3786 5216 3792 5228
rect 3467 5188 3792 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 5000 5216 5028 5324
rect 5445 5321 5457 5324
rect 5491 5352 5503 5355
rect 7190 5352 7196 5364
rect 5491 5324 7196 5352
rect 5491 5321 5503 5324
rect 5445 5315 5503 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8386 5352 8392 5364
rect 8067 5324 8392 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 6730 5284 6736 5296
rect 5736 5256 6736 5284
rect 4816 5188 5028 5216
rect 5169 5219 5227 5225
rect 4816 5160 4844 5188
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5442 5216 5448 5228
rect 5215 5188 5448 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 4798 5108 4804 5160
rect 4856 5108 4862 5160
rect 5736 5157 5764 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 6825 5287 6883 5293
rect 6825 5253 6837 5287
rect 6871 5253 6883 5287
rect 6825 5247 6883 5253
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5148 6699 5151
rect 6840 5148 6868 5247
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 8036 5216 8064 5315
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 8904 5324 10364 5352
rect 8904 5312 8910 5324
rect 8110 5244 8116 5296
rect 8168 5244 8174 5296
rect 10336 5284 10364 5324
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10468 5324 10517 5352
rect 10468 5312 10474 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 12526 5352 12532 5364
rect 10505 5315 10563 5321
rect 11440 5324 12532 5352
rect 10594 5284 10600 5296
rect 10336 5256 10600 5284
rect 10594 5244 10600 5256
rect 10652 5244 10658 5296
rect 7515 5188 8064 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 6687 5120 6868 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6972 5120 7205 5148
rect 6972 5108 6978 5120
rect 7193 5117 7205 5120
rect 7239 5148 7251 5151
rect 8128 5148 8156 5244
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9398 5216 9404 5228
rect 8803 5188 9404 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9398 5176 9404 5188
rect 9456 5216 9462 5228
rect 9674 5216 9680 5228
rect 9456 5188 9680 5216
rect 9456 5176 9462 5188
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10836 5188 10977 5216
rect 10836 5176 10842 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 7239 5120 8156 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10744 5120 10885 5148
rect 10744 5108 10750 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 7285 5083 7343 5089
rect 7285 5049 7297 5083
rect 7331 5080 7343 5083
rect 8018 5080 8024 5092
rect 7331 5052 8024 5080
rect 7331 5049 7343 5052
rect 7285 5043 7343 5049
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8113 5083 8171 5089
rect 8113 5049 8125 5083
rect 8159 5049 8171 5083
rect 8113 5043 8171 5049
rect 9033 5083 9091 5089
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9306 5080 9312 5092
rect 9079 5052 9312 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 8128 5012 8156 5043
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9490 5040 9496 5092
rect 9548 5040 9554 5092
rect 10888 5080 10916 5111
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 11112 5120 11161 5148
rect 11112 5108 11118 5120
rect 11149 5117 11161 5120
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 11440 5089 11468 5324
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13412 5324 15884 5352
rect 13412 5312 13418 5324
rect 15856 5296 15884 5324
rect 16114 5312 16120 5364
rect 16172 5312 16178 5364
rect 16853 5355 16911 5361
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 18414 5352 18420 5364
rect 16899 5324 18420 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 18414 5312 18420 5324
rect 18472 5312 18478 5364
rect 11606 5244 11612 5296
rect 11664 5244 11670 5296
rect 11701 5287 11759 5293
rect 11701 5253 11713 5287
rect 11747 5284 11759 5287
rect 13814 5284 13820 5296
rect 11747 5256 13820 5284
rect 11747 5253 11759 5256
rect 11701 5247 11759 5253
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 14090 5244 14096 5296
rect 14148 5284 14154 5296
rect 15654 5284 15660 5296
rect 14148 5256 15660 5284
rect 14148 5244 14154 5256
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 15746 5244 15752 5296
rect 15804 5244 15810 5296
rect 15838 5244 15844 5296
rect 15896 5284 15902 5296
rect 16206 5284 16212 5296
rect 15896 5256 16212 5284
rect 15896 5244 15902 5256
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 11624 5157 11652 5244
rect 11716 5188 11836 5216
rect 11716 5157 11744 5188
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5117 11667 5151
rect 11609 5111 11667 5117
rect 11701 5151 11759 5157
rect 11701 5117 11713 5151
rect 11747 5117 11759 5151
rect 11808 5148 11836 5188
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 16393 5219 16451 5225
rect 12768 5188 15976 5216
rect 12768 5176 12774 5188
rect 11974 5148 11980 5160
rect 11808 5120 11980 5148
rect 11701 5111 11759 5117
rect 11425 5083 11483 5089
rect 11425 5080 11437 5083
rect 10888 5052 11437 5080
rect 11425 5049 11437 5052
rect 11471 5049 11483 5083
rect 11624 5080 11652 5111
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 12250 5108 12256 5160
rect 12308 5108 12314 5160
rect 12986 5148 12992 5160
rect 12406 5120 12992 5148
rect 12406 5080 12434 5120
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 14277 5151 14335 5157
rect 13403 5120 13676 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 11624 5052 12434 5080
rect 11425 5043 11483 5049
rect 9398 5012 9404 5024
rect 8128 4984 9404 5012
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 11330 4972 11336 5024
rect 11388 4972 11394 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11974 5012 11980 5024
rect 11572 4984 11980 5012
rect 11572 4972 11578 4984
rect 11974 4972 11980 4984
rect 12032 5012 12038 5024
rect 12986 5012 12992 5024
rect 12032 4984 12992 5012
rect 12032 4972 12038 4984
rect 12986 4972 12992 4984
rect 13044 5012 13050 5024
rect 13354 5012 13360 5024
rect 13044 4984 13360 5012
rect 13044 4972 13050 4984
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13648 5021 13676 5120
rect 14277 5117 14289 5151
rect 14323 5148 14335 5151
rect 15286 5148 15292 5160
rect 14323 5120 15292 5148
rect 14323 5117 14335 5120
rect 14277 5111 14335 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15378 5108 15384 5160
rect 15436 5108 15442 5160
rect 15948 5157 15976 5188
rect 16393 5185 16405 5219
rect 16439 5185 16451 5219
rect 16393 5179 16451 5185
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5216 18475 5219
rect 18463 5188 18552 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 16298 5108 16304 5160
rect 16356 5108 16362 5160
rect 13909 5083 13967 5089
rect 13909 5049 13921 5083
rect 13955 5080 13967 5083
rect 13998 5080 14004 5092
rect 13955 5052 14004 5080
rect 13955 5049 13967 5052
rect 13909 5043 13967 5049
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 15654 5040 15660 5092
rect 15712 5080 15718 5092
rect 16408 5080 16436 5179
rect 18524 5160 18552 5188
rect 16574 5108 16580 5160
rect 16632 5108 16638 5160
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5148 17003 5151
rect 17494 5148 17500 5160
rect 16991 5120 17500 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 16482 5080 16488 5092
rect 15712 5052 16488 5080
rect 15712 5040 15718 5052
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 16684 5080 16712 5111
rect 17494 5108 17500 5120
rect 17552 5108 17558 5160
rect 17586 5108 17592 5160
rect 17644 5108 17650 5160
rect 18506 5108 18512 5160
rect 18564 5108 18570 5160
rect 18782 5108 18788 5160
rect 18840 5108 18846 5160
rect 18966 5108 18972 5160
rect 19024 5108 19030 5160
rect 17402 5080 17408 5092
rect 16684 5052 17408 5080
rect 17402 5040 17408 5052
rect 17460 5040 17466 5092
rect 17604 5080 17632 5108
rect 18046 5080 18052 5092
rect 17604 5052 18052 5080
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 18693 5083 18751 5089
rect 18693 5049 18705 5083
rect 18739 5049 18751 5083
rect 18693 5043 18751 5049
rect 13633 5015 13691 5021
rect 13633 4981 13645 5015
rect 13679 5012 13691 5015
rect 14274 5012 14280 5024
rect 13679 4984 14280 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 18708 5012 18736 5043
rect 17276 4984 18736 5012
rect 17276 4972 17282 4984
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 6454 4808 6460 4820
rect 3844 4780 6040 4808
rect 3844 4768 3850 4780
rect 474 4632 480 4684
rect 532 4672 538 4684
rect 3896 4681 3924 4780
rect 4157 4743 4215 4749
rect 4157 4709 4169 4743
rect 4203 4740 4215 4743
rect 4430 4740 4436 4752
rect 4203 4712 4436 4740
rect 4203 4709 4215 4712
rect 4157 4703 4215 4709
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 4798 4700 4804 4752
rect 4856 4700 4862 4752
rect 6012 4681 6040 4780
rect 6288 4780 6460 4808
rect 6288 4749 6316 4780
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7745 4811 7803 4817
rect 7248 4780 7420 4808
rect 7248 4768 7254 4780
rect 6273 4743 6331 4749
rect 6273 4709 6285 4743
rect 6319 4709 6331 4743
rect 6273 4703 6331 4709
rect 845 4675 903 4681
rect 845 4672 857 4675
rect 532 4644 857 4672
rect 532 4632 538 4644
rect 845 4641 857 4644
rect 891 4641 903 4675
rect 845 4635 903 4641
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4641 3939 4675
rect 3881 4635 3939 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 7392 4658 7420 4780
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8018 4808 8024 4820
rect 7791 4780 8024 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 10410 4808 10416 4820
rect 8987 4780 10416 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 11422 4808 11428 4820
rect 10827 4780 11428 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11698 4768 11704 4820
rect 11756 4768 11762 4820
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 12250 4808 12256 4820
rect 11848 4780 12256 4808
rect 11848 4768 11854 4780
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 16114 4768 16120 4820
rect 16172 4768 16178 4820
rect 16206 4768 16212 4820
rect 16264 4768 16270 4820
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 17862 4808 17868 4820
rect 17460 4780 17868 4808
rect 17460 4768 17466 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 10962 4740 10968 4752
rect 8220 4712 10968 4740
rect 8220 4681 8248 4712
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11057 4743 11115 4749
rect 11057 4709 11069 4743
rect 11103 4740 11115 4743
rect 12069 4743 12127 4749
rect 12069 4740 12081 4743
rect 11103 4712 12081 4740
rect 11103 4709 11115 4712
rect 11057 4703 11115 4709
rect 12069 4709 12081 4712
rect 12115 4709 12127 4743
rect 12069 4703 12127 4709
rect 12158 4700 12164 4752
rect 12216 4740 12222 4752
rect 16132 4740 16160 4768
rect 12216 4712 12558 4740
rect 15856 4712 16160 4740
rect 12216 4700 12222 4712
rect 8205 4675 8263 4681
rect 5997 4635 6055 4641
rect 8205 4641 8217 4675
rect 8251 4641 8263 4675
rect 8205 4635 8263 4641
rect 8294 4632 8300 4684
rect 8352 4632 8358 4684
rect 9668 4675 9726 4681
rect 8772 4644 9260 4672
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 7926 4604 7932 4616
rect 5675 4576 7932 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8772 4613 8800 4644
rect 9232 4616 9260 4644
rect 9668 4641 9680 4675
rect 9714 4672 9726 4675
rect 10226 4672 10232 4684
rect 9714 4644 10232 4672
rect 9714 4641 9726 4644
rect 9668 4635 9726 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 11606 4672 11612 4684
rect 11379 4644 11612 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15378 4672 15384 4684
rect 14783 4644 15384 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 15856 4681 15884 4712
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 16724 4712 17540 4740
rect 16724 4700 16730 4712
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 15930 4632 15936 4684
rect 15988 4672 15994 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15988 4644 16129 4672
rect 15988 4632 15994 4644
rect 16117 4641 16129 4644
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16356 4644 16405 4672
rect 16356 4632 16362 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 16899 4644 17080 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 8846 4564 8852 4616
rect 8904 4564 8910 4616
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9398 4564 9404 4616
rect 9456 4564 9462 4616
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11112 4576 11253 4604
rect 11112 4564 11118 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 12526 4604 12532 4616
rect 11839 4576 12532 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 13780 4576 13829 4604
rect 13780 4564 13786 4576
rect 13817 4573 13829 4576
rect 13863 4604 13875 4607
rect 15948 4604 15976 4632
rect 13863 4576 15976 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 16482 4564 16488 4616
rect 16540 4604 16546 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16540 4576 16957 4604
rect 16540 4564 16546 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 17052 4604 17080 4644
rect 17126 4632 17132 4684
rect 17184 4632 17190 4684
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4672 17279 4675
rect 17310 4672 17316 4684
rect 17267 4644 17316 4672
rect 17267 4641 17279 4644
rect 17221 4635 17279 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17512 4681 17540 4712
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4641 17555 4675
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 17497 4635 17555 4641
rect 17926 4644 19073 4672
rect 17926 4604 17954 4644
rect 19061 4641 19073 4644
rect 19107 4672 19119 4675
rect 19150 4672 19156 4684
rect 19107 4644 19156 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 17052 4576 17954 4604
rect 16945 4567 17003 4573
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18506 4604 18512 4616
rect 18104 4576 18512 4604
rect 18104 4564 18110 4576
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 14553 4539 14611 4545
rect 14553 4505 14565 4539
rect 14599 4536 14611 4539
rect 14826 4536 14832 4548
rect 14599 4508 14832 4536
rect 14599 4505 14611 4508
rect 14553 4499 14611 4505
rect 14826 4496 14832 4508
rect 14884 4496 14890 4548
rect 1026 4428 1032 4480
rect 1084 4428 1090 4480
rect 8478 4428 8484 4480
rect 8536 4428 8542 4480
rect 9309 4471 9367 4477
rect 9309 4437 9321 4471
rect 9355 4468 9367 4471
rect 10410 4468 10416 4480
rect 9355 4440 10416 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 11146 4468 11152 4480
rect 10560 4440 11152 4468
rect 10560 4428 10566 4440
rect 11146 4428 11152 4440
rect 11204 4468 11210 4480
rect 12158 4468 12164 4480
rect 11204 4440 12164 4468
rect 11204 4428 11210 4440
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 14918 4428 14924 4480
rect 14976 4468 14982 4480
rect 16577 4471 16635 4477
rect 16577 4468 16589 4471
rect 14976 4440 16589 4468
rect 14976 4428 14982 4440
rect 16577 4437 16589 4440
rect 16623 4437 16635 4471
rect 16577 4431 16635 4437
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 12802 4264 12808 4276
rect 8352 4236 12808 4264
rect 8352 4224 8358 4236
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 17770 4224 17776 4276
rect 17828 4264 17834 4276
rect 18233 4267 18291 4273
rect 18233 4264 18245 4267
rect 17828 4236 18245 4264
rect 17828 4224 17834 4236
rect 18233 4233 18245 4236
rect 18279 4233 18291 4267
rect 18233 4227 18291 4233
rect 9214 4156 9220 4208
rect 9272 4196 9278 4208
rect 9309 4199 9367 4205
rect 9309 4196 9321 4199
rect 9272 4168 9321 4196
rect 9272 4156 9278 4168
rect 9309 4165 9321 4168
rect 9355 4165 9367 4199
rect 10686 4196 10692 4208
rect 9309 4159 9367 4165
rect 9876 4168 10692 4196
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 6273 4131 6331 4137
rect 900 4100 1532 4128
rect 900 4088 906 4100
rect 1026 4020 1032 4072
rect 1084 4020 1090 4072
rect 1136 4069 1164 4100
rect 1121 4063 1179 4069
rect 1121 4029 1133 4063
rect 1167 4029 1179 4063
rect 1121 4023 1179 4029
rect 1213 4063 1271 4069
rect 1213 4029 1225 4063
rect 1259 4060 1271 4063
rect 1397 4063 1455 4069
rect 1397 4060 1409 4063
rect 1259 4032 1409 4060
rect 1259 4029 1271 4032
rect 1213 4023 1271 4029
rect 1397 4029 1409 4032
rect 1443 4029 1455 4063
rect 1504 4060 1532 4100
rect 2792 4100 3372 4128
rect 2792 4060 2820 4100
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 1504 4032 2881 4060
rect 1397 4023 1455 4029
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4060 3019 4063
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3007 4032 3249 4060
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 3344 4060 3372 4100
rect 6273 4097 6285 4131
rect 6319 4128 6331 4131
rect 7282 4128 7288 4140
rect 6319 4100 7288 4128
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8202 4128 8208 4140
rect 8067 4100 8208 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 8260 4100 8861 4128
rect 8260 4088 8266 4100
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9079 4100 9628 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9600 4072 9628 4100
rect 3786 4060 3792 4072
rect 3344 4032 3792 4060
rect 3237 4023 3295 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 7984 4032 8769 4060
rect 7984 4020 7990 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 9582 4020 9588 4072
rect 9640 4020 9646 4072
rect 9876 4069 9904 4168
rect 10686 4156 10692 4168
rect 10744 4196 10750 4208
rect 10744 4168 12434 4196
rect 10744 4156 10750 4168
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4128 10011 4131
rect 11054 4128 11060 4140
rect 9999 4100 11060 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4128 11667 4131
rect 11974 4128 11980 4140
rect 11655 4100 11980 4128
rect 11655 4097 11667 4100
rect 11609 4091 11667 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10226 4060 10232 4072
rect 10183 4032 10232 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 1044 3992 1072 4020
rect 1642 3995 1700 4001
rect 1642 3992 1654 3995
rect 1044 3964 1654 3992
rect 1642 3961 1654 3964
rect 1688 3961 1700 3995
rect 1642 3955 1700 3961
rect 3504 3995 3562 4001
rect 3504 3961 3516 3995
rect 3550 3992 3562 3995
rect 3602 3992 3608 4004
rect 3550 3964 3608 3992
rect 3550 3961 3562 3964
rect 3504 3955 3562 3961
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 6546 3952 6552 4004
rect 6604 3952 6610 4004
rect 7190 3952 7196 4004
rect 7248 3952 7254 4004
rect 10060 3992 10088 4023
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 11532 3992 11560 4088
rect 11698 4020 11704 4072
rect 11756 4020 11762 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 10060 3964 11560 3992
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 4890 3924 4896 3936
rect 4663 3896 4896 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8168 3896 8401 3924
rect 8168 3884 8174 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 10502 3924 10508 3936
rect 9272 3896 10508 3924
rect 9272 3884 9278 3896
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11808 3924 11836 4023
rect 12406 3992 12434 4168
rect 12618 4156 12624 4208
rect 12676 4156 12682 4208
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 15381 4199 15439 4205
rect 15381 4196 15393 4199
rect 14884 4168 15393 4196
rect 14884 4156 14890 4168
rect 15381 4165 15393 4168
rect 15427 4196 15439 4199
rect 16666 4196 16672 4208
rect 15427 4168 16672 4196
rect 15427 4165 15439 4168
rect 15381 4159 15439 4165
rect 12636 4060 12664 4156
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13998 4128 14004 4140
rect 13403 4100 14004 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13722 4060 13728 4072
rect 12636 4032 13728 4060
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 12406 3964 13645 3992
rect 13633 3961 13645 3964
rect 13679 3961 13691 3995
rect 13633 3955 13691 3961
rect 11572 3896 11836 3924
rect 13832 3924 13860 4100
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 15488 4069 15516 4168
rect 16666 4156 16672 4168
rect 16724 4196 16730 4208
rect 17037 4199 17095 4205
rect 17037 4196 17049 4199
rect 16724 4168 17049 4196
rect 16724 4156 16730 4168
rect 17037 4165 17049 4168
rect 17083 4196 17095 4199
rect 18046 4196 18052 4208
rect 17083 4168 18052 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4128 15623 4131
rect 15611 4100 16804 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 13924 3992 13952 4023
rect 15580 3992 15608 4091
rect 16666 4020 16672 4072
rect 16724 4020 16730 4072
rect 16776 4060 16804 4100
rect 17218 4060 17224 4072
rect 16776 4032 17224 4060
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 18690 4060 18696 4072
rect 18463 4032 18696 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 18874 4020 18880 4072
rect 18932 4020 18938 4072
rect 13924 3964 15608 3992
rect 16206 3952 16212 4004
rect 16264 3992 16270 4004
rect 17313 3995 17371 4001
rect 17313 3992 17325 3995
rect 16264 3964 17325 3992
rect 16264 3952 16270 3964
rect 17313 3961 17325 3964
rect 17359 3961 17371 3995
rect 18141 3995 18199 4001
rect 18141 3992 18153 3995
rect 17313 3955 17371 3961
rect 17926 3964 18153 3992
rect 17926 3924 17954 3964
rect 18141 3961 18153 3964
rect 18187 3992 18199 3995
rect 18187 3964 18828 3992
rect 18187 3961 18199 3964
rect 18141 3955 18199 3961
rect 18800 3933 18828 3964
rect 13832 3896 17954 3924
rect 18785 3927 18843 3933
rect 11572 3884 11578 3896
rect 18785 3893 18797 3927
rect 18831 3893 18843 3927
rect 18785 3887 18843 3893
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 2774 3680 2780 3732
rect 2832 3680 2838 3732
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3660 3692 3801 3720
rect 3660 3680 3666 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 3789 3683 3847 3689
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 6604 3692 6745 3720
rect 6604 3680 6610 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 6733 3683 6791 3689
rect 8110 3680 8116 3732
rect 8168 3680 8174 3732
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11204 3692 12572 3720
rect 11204 3680 11210 3692
rect 2792 3584 2820 3680
rect 3145 3587 3203 3593
rect 3145 3584 3157 3587
rect 2792 3556 3157 3584
rect 3145 3553 3157 3556
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 8128 3584 8156 3680
rect 8570 3612 8576 3664
rect 8628 3612 8634 3664
rect 9692 3652 9720 3680
rect 10502 3652 10508 3664
rect 9692 3624 9904 3652
rect 9876 3593 9904 3624
rect 10336 3624 10508 3652
rect 10336 3593 10364 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 11241 3655 11299 3661
rect 11241 3621 11253 3655
rect 11287 3652 11299 3655
rect 11330 3652 11336 3664
rect 11287 3624 11336 3652
rect 11287 3621 11299 3624
rect 11241 3615 11299 3621
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 12544 3652 12572 3692
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 15841 3723 15899 3729
rect 13780 3692 15148 3720
rect 13780 3680 13786 3692
rect 12466 3624 13846 3652
rect 14918 3612 14924 3664
rect 14976 3612 14982 3664
rect 15120 3661 15148 3692
rect 15841 3689 15853 3723
rect 15887 3720 15899 3723
rect 16298 3720 16304 3732
rect 15887 3692 16304 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 17494 3680 17500 3732
rect 17552 3680 17558 3732
rect 15105 3655 15163 3661
rect 15105 3621 15117 3655
rect 15151 3621 15163 3655
rect 15105 3615 15163 3621
rect 6963 3556 8156 3584
rect 9861 3587 9919 3593
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 9861 3553 9873 3587
rect 9907 3584 9919 3587
rect 10137 3587 10195 3593
rect 9907 3556 10088 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8846 3516 8852 3528
rect 8159 3488 8852 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 9631 3488 9996 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 9968 3457 9996 3488
rect 9953 3451 10011 3457
rect 9953 3417 9965 3451
rect 9999 3417 10011 3451
rect 10060 3448 10088 3556
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 10152 3516 10180 3547
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10520 3556 10977 3584
rect 10428 3516 10456 3544
rect 10152 3488 10456 3516
rect 10520 3448 10548 3556
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 10965 3547 11023 3553
rect 12544 3556 13093 3584
rect 10980 3516 11008 3547
rect 12544 3528 12572 3556
rect 13081 3553 13093 3556
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 12526 3516 12532 3528
rect 10980 3488 12532 3516
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12986 3476 12992 3528
rect 13044 3476 13050 3528
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14936 3516 14964 3612
rect 15120 3584 15148 3615
rect 15197 3587 15255 3593
rect 15197 3584 15209 3587
rect 15120 3556 15209 3584
rect 15197 3553 15209 3556
rect 15243 3553 15255 3587
rect 15197 3547 15255 3553
rect 17402 3544 17408 3596
rect 17460 3544 17466 3596
rect 17586 3544 17592 3596
rect 17644 3544 17650 3596
rect 18138 3544 18144 3596
rect 18196 3584 18202 3596
rect 18509 3587 18567 3593
rect 18509 3584 18521 3587
rect 18196 3556 18521 3584
rect 18196 3544 18202 3556
rect 18509 3553 18521 3556
rect 18555 3553 18567 3587
rect 18509 3547 18567 3553
rect 18598 3544 18604 3596
rect 18656 3544 18662 3596
rect 13403 3488 14964 3516
rect 17957 3519 18015 3525
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 18003 3488 18245 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18233 3485 18245 3488
rect 18279 3516 18291 3519
rect 18616 3516 18644 3544
rect 18279 3488 18644 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 10060 3420 10548 3448
rect 9953 3411 10011 3417
rect 10778 3408 10784 3460
rect 10836 3408 10842 3460
rect 10597 3383 10655 3389
rect 10597 3349 10609 3383
rect 10643 3380 10655 3383
rect 13004 3380 13032 3476
rect 10643 3352 13032 3380
rect 10643 3349 10655 3352
rect 10597 3343 10655 3349
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 16206 3176 16212 3188
rect 14936 3148 16212 3176
rect 7392 3040 7420 3136
rect 14936 3120 14964 3148
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 16758 3136 16764 3188
rect 16816 3136 16822 3188
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 14918 3108 14924 3120
rect 7892 3080 14924 3108
rect 7892 3068 7898 3080
rect 8496 3049 8524 3080
rect 8481 3043 8539 3049
rect 7392 3012 8248 3040
rect 8220 2984 8248 3012
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3040 10195 3043
rect 10226 3040 10232 3052
rect 10183 3012 10232 3040
rect 10183 3009 10195 3012
rect 10137 3003 10195 3009
rect 6822 2932 6828 2984
rect 6880 2932 6886 2984
rect 7006 2932 7012 2984
rect 7064 2932 7070 2984
rect 7282 2932 7288 2984
rect 7340 2932 7346 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 7576 2904 7604 2935
rect 8202 2932 8208 2984
rect 8260 2932 8266 2984
rect 7248 2876 7604 2904
rect 9968 2904 9996 3003
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11422 3000 11428 3052
rect 11480 3000 11486 3052
rect 11809 3049 11837 3080
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 15120 3080 16344 3108
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 15120 3049 15148 3080
rect 13265 3043 13323 3049
rect 13265 3040 13277 3043
rect 12032 3012 13277 3040
rect 12032 3000 12038 3012
rect 13265 3009 13277 3012
rect 13311 3040 13323 3043
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13311 3012 13921 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 15105 3043 15163 3049
rect 15105 3009 15117 3043
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 16206 3040 16212 3052
rect 15795 3012 16212 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 10045 2975 10103 2981
rect 10045 2941 10057 2975
rect 10091 2972 10103 2975
rect 11514 2972 11520 2984
rect 10091 2944 11520 2972
rect 10091 2941 10103 2944
rect 10045 2935 10103 2941
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11609 2975 11667 2981
rect 11609 2941 11621 2975
rect 11655 2941 11667 2975
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 11609 2935 11667 2941
rect 12820 2944 12909 2972
rect 10686 2904 10692 2916
rect 9968 2876 10692 2904
rect 7248 2864 7254 2876
rect 10686 2864 10692 2876
rect 10744 2864 10750 2916
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 7800 2808 8125 2836
rect 7800 2796 7806 2808
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 11532 2836 11560 2932
rect 11624 2904 11652 2935
rect 11698 2904 11704 2916
rect 11624 2876 11704 2904
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 12820 2904 12848 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 13924 2972 13952 3003
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13924 2944 14013 2972
rect 12897 2935 12955 2941
rect 14001 2941 14013 2944
rect 14047 2972 14059 2975
rect 14090 2972 14096 2984
rect 14047 2944 14096 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14090 2932 14096 2944
rect 14148 2972 14154 2984
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 14148 2944 15669 2972
rect 14148 2932 14154 2944
rect 15657 2941 15669 2944
rect 15703 2972 15715 2975
rect 15764 2972 15792 3003
rect 16206 3000 16212 3012
rect 16264 3000 16270 3052
rect 15703 2944 15792 2972
rect 16316 2972 16344 3080
rect 16776 3040 16804 3136
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16776 3012 16865 3040
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17218 3000 17224 3052
rect 17276 3000 17282 3052
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 16316 2944 16773 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16761 2941 16773 2944
rect 16807 2972 16819 2975
rect 17236 2972 17264 3000
rect 16807 2944 17264 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 17954 2932 17960 2984
rect 18012 2932 18018 2984
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2972 19119 2975
rect 19702 2972 19708 2984
rect 19107 2944 19708 2972
rect 19107 2941 19119 2944
rect 19061 2935 19119 2941
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 14458 2904 14464 2916
rect 12820 2876 14464 2904
rect 12820 2836 12848 2876
rect 14458 2864 14464 2876
rect 14516 2904 14522 2916
rect 17494 2904 17500 2916
rect 14516 2876 17500 2904
rect 14516 2864 14522 2876
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 11532 2808 12848 2836
rect 8113 2799 8171 2805
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 18877 2839 18935 2845
rect 18877 2836 18889 2839
rect 13964 2808 18889 2836
rect 13964 2796 13970 2808
rect 18877 2805 18889 2808
rect 18923 2805 18935 2839
rect 18877 2799 18935 2805
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 18877 2635 18935 2641
rect 18877 2632 18889 2635
rect 16632 2604 18889 2632
rect 16632 2592 16638 2604
rect 18877 2601 18889 2604
rect 18923 2601 18935 2635
rect 18877 2595 18935 2601
rect 6730 2564 6736 2576
rect 5828 2536 6736 2564
rect 5828 2505 5856 2536
rect 6104 2508 6132 2536
rect 6730 2524 6736 2536
rect 6788 2524 6794 2576
rect 6822 2524 6828 2576
rect 6880 2564 6886 2576
rect 7990 2567 8048 2573
rect 7990 2564 8002 2567
rect 6880 2536 8002 2564
rect 6880 2524 6886 2536
rect 7990 2533 8002 2536
rect 8036 2533 8048 2567
rect 7990 2527 8048 2533
rect 12406 2536 14412 2564
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 6012 2428 6040 2459
rect 6086 2456 6092 2508
rect 6144 2456 6150 2508
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2496 6331 2499
rect 6641 2499 6699 2505
rect 6641 2496 6653 2499
rect 6319 2468 6653 2496
rect 6319 2465 6331 2468
rect 6273 2459 6331 2465
rect 6641 2465 6653 2468
rect 6687 2465 6699 2499
rect 6641 2459 6699 2465
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 7064 2468 7205 2496
rect 7064 2456 7070 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 7742 2456 7748 2508
rect 7800 2456 7806 2508
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 10318 2496 10324 2508
rect 9263 2468 10324 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 10827 2468 11437 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 11425 2465 11437 2468
rect 11471 2496 11483 2499
rect 12406 2496 12434 2536
rect 11471 2468 12434 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 13170 2496 13176 2508
rect 12676 2468 13176 2496
rect 12676 2456 12682 2468
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 14090 2456 14096 2508
rect 14148 2456 14154 2508
rect 14384 2505 14412 2536
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 15838 2496 15844 2508
rect 14415 2468 15844 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 15838 2456 15844 2468
rect 15896 2496 15902 2508
rect 17221 2499 17279 2505
rect 17221 2496 17233 2499
rect 15896 2468 17233 2496
rect 15896 2456 15902 2468
rect 17221 2465 17233 2468
rect 17267 2465 17279 2499
rect 17221 2459 17279 2465
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 6012 2400 7481 2428
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10686 2428 10692 2440
rect 10643 2400 10692 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10686 2388 10692 2400
rect 10744 2428 10750 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10744 2400 11529 2428
rect 10744 2388 10750 2400
rect 11517 2397 11529 2400
rect 11563 2428 11575 2431
rect 11606 2428 11612 2440
rect 11563 2400 11612 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11974 2388 11980 2440
rect 12032 2428 12038 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12032 2400 12541 2428
rect 12032 2388 12038 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 14001 2431 14059 2437
rect 14001 2397 14013 2431
rect 14047 2428 14059 2431
rect 14108 2428 14136 2456
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14047 2400 14565 2428
rect 14047 2397 14059 2400
rect 14001 2391 14059 2397
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 15746 2428 15752 2440
rect 14553 2391 14611 2397
rect 15166 2400 15752 2428
rect 12544 2360 12572 2391
rect 14458 2360 14464 2372
rect 12544 2332 14464 2360
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 6914 2252 6920 2304
rect 6972 2252 6978 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 11514 2292 11520 2304
rect 9171 2264 11520 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 14476 2292 14504 2320
rect 15166 2292 15194 2400
rect 15746 2388 15752 2400
rect 15804 2428 15810 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15804 2400 15945 2428
rect 15804 2388 15810 2400
rect 15933 2397 15945 2400
rect 15979 2428 15991 2431
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15979 2400 16129 2428
rect 15979 2397 15991 2400
rect 15933 2391 15991 2397
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 17236 2428 17264 2459
rect 18322 2456 18328 2508
rect 18380 2456 18386 2508
rect 19061 2499 19119 2505
rect 19061 2465 19073 2499
rect 19107 2496 19119 2499
rect 19610 2496 19616 2508
rect 19107 2468 19616 2496
rect 19107 2465 19119 2468
rect 19061 2459 19119 2465
rect 19610 2456 19616 2468
rect 19668 2456 19674 2508
rect 18230 2428 18236 2440
rect 17236 2400 18236 2428
rect 16117 2391 16175 2397
rect 18230 2388 18236 2400
rect 18288 2428 18294 2440
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18288 2400 18521 2428
rect 18288 2388 18294 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 17589 2363 17647 2369
rect 17589 2329 17601 2363
rect 17635 2360 17647 2363
rect 17862 2360 17868 2372
rect 17635 2332 17868 2360
rect 17635 2329 17647 2332
rect 17589 2323 17647 2329
rect 17862 2320 17868 2332
rect 17920 2320 17926 2372
rect 14476 2264 15194 2292
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 6503 2091 6561 2097
rect 6503 2057 6515 2091
rect 6549 2088 6561 2091
rect 6822 2088 6828 2100
rect 6549 2060 6828 2088
rect 6549 2057 6561 2060
rect 6503 2051 6561 2057
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 6914 2048 6920 2100
rect 6972 2048 6978 2100
rect 8113 2091 8171 2097
rect 8113 2057 8125 2091
rect 8159 2088 8171 2091
rect 9398 2088 9404 2100
rect 8159 2060 9404 2088
rect 8159 2057 8171 2060
rect 8113 2051 8171 2057
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 11790 2088 11796 2100
rect 10152 2060 11796 2088
rect 6932 2020 6960 2048
rect 10152 2020 10180 2060
rect 11790 2048 11796 2060
rect 11848 2088 11854 2100
rect 15010 2088 15016 2100
rect 11848 2060 15016 2088
rect 11848 2048 11854 2060
rect 15010 2048 15016 2060
rect 15068 2048 15074 2100
rect 6288 1992 6960 2020
rect 8680 1992 10180 2020
rect 14001 2023 14059 2029
rect 842 1844 848 1896
rect 900 1844 906 1896
rect 5718 1844 5724 1896
rect 5776 1844 5782 1896
rect 5810 1844 5816 1896
rect 5868 1844 5874 1896
rect 6288 1893 6316 1992
rect 6963 1955 7021 1961
rect 6963 1952 6975 1955
rect 6656 1924 6975 1952
rect 6089 1887 6147 1893
rect 6089 1853 6101 1887
rect 6135 1853 6147 1887
rect 6089 1847 6147 1853
rect 6273 1887 6331 1893
rect 6273 1853 6285 1887
rect 6319 1853 6331 1887
rect 6273 1847 6331 1853
rect 6432 1887 6490 1893
rect 6432 1853 6444 1887
rect 6478 1884 6490 1887
rect 6656 1884 6684 1924
rect 6963 1921 6975 1924
rect 7009 1921 7021 1955
rect 6963 1915 7021 1921
rect 8680 1896 8708 1992
rect 14001 1989 14013 2023
rect 14047 2020 14059 2023
rect 14182 2020 14188 2032
rect 14047 1992 14188 2020
rect 14047 1989 14059 1992
rect 14001 1983 14059 1989
rect 14182 1980 14188 1992
rect 14240 1980 14246 2032
rect 16206 1980 16212 2032
rect 16264 2020 16270 2032
rect 17862 2020 17868 2032
rect 16264 1992 17868 2020
rect 16264 1980 16270 1992
rect 17862 1980 17868 1992
rect 17920 2020 17926 2032
rect 17920 1992 18092 2020
rect 17920 1980 17926 1992
rect 8849 1955 8907 1961
rect 8849 1921 8861 1955
rect 8895 1921 8907 1955
rect 8849 1915 8907 1921
rect 6478 1856 6684 1884
rect 6825 1887 6883 1893
rect 6478 1853 6490 1856
rect 6432 1847 6490 1853
rect 6825 1853 6837 1887
rect 6871 1853 6883 1887
rect 6825 1847 6883 1853
rect 7066 1887 7124 1893
rect 7066 1853 7078 1887
rect 7112 1884 7124 1887
rect 7282 1884 7288 1896
rect 7112 1856 7288 1884
rect 7112 1853 7124 1856
rect 7066 1847 7124 1853
rect 6104 1760 6132 1847
rect 6840 1816 6868 1847
rect 7282 1844 7288 1856
rect 7340 1844 7346 1896
rect 7374 1844 7380 1896
rect 7432 1844 7438 1896
rect 7466 1844 7472 1896
rect 7524 1844 7530 1896
rect 7926 1844 7932 1896
rect 7984 1844 7990 1896
rect 8018 1844 8024 1896
rect 8076 1844 8082 1896
rect 8662 1844 8668 1896
rect 8720 1844 8726 1896
rect 8864 1884 8892 1915
rect 11606 1912 11612 1964
rect 11664 1952 11670 1964
rect 13265 1955 13323 1961
rect 13265 1952 13277 1955
rect 11664 1924 13277 1952
rect 11664 1912 11670 1924
rect 8941 1887 8999 1893
rect 8941 1884 8953 1887
rect 8864 1856 8953 1884
rect 8941 1853 8953 1856
rect 8987 1884 8999 1887
rect 9030 1884 9036 1896
rect 8987 1856 9036 1884
rect 8987 1853 8999 1856
rect 8941 1847 8999 1853
rect 9030 1844 9036 1856
rect 9088 1844 9094 1896
rect 9674 1844 9680 1896
rect 9732 1884 9738 1896
rect 10045 1887 10103 1893
rect 10045 1884 10057 1887
rect 9732 1856 10057 1884
rect 9732 1844 9738 1856
rect 10045 1853 10057 1856
rect 10091 1884 10103 1887
rect 10137 1887 10195 1893
rect 10137 1884 10149 1887
rect 10091 1856 10149 1884
rect 10091 1853 10103 1856
rect 10045 1847 10103 1853
rect 10137 1853 10149 1856
rect 10183 1884 10195 1887
rect 10870 1884 10876 1896
rect 10183 1856 10876 1884
rect 10183 1853 10195 1856
rect 10137 1847 10195 1853
rect 10870 1844 10876 1856
rect 10928 1844 10934 1896
rect 11716 1893 11744 1924
rect 13265 1921 13277 1924
rect 13311 1952 13323 1955
rect 13630 1952 13636 1964
rect 13311 1924 13636 1952
rect 13311 1921 13323 1924
rect 13265 1915 13323 1921
rect 13630 1912 13636 1924
rect 13688 1952 13694 1964
rect 14090 1952 14096 1964
rect 13688 1924 14096 1952
rect 13688 1912 13694 1924
rect 14090 1912 14096 1924
rect 14148 1912 14154 1964
rect 16758 1912 16764 1964
rect 16816 1952 16822 1964
rect 18064 1961 18092 1992
rect 16853 1955 16911 1961
rect 16853 1952 16865 1955
rect 16816 1924 16865 1952
rect 16816 1912 16822 1924
rect 16853 1921 16865 1924
rect 16899 1921 16911 1955
rect 16853 1915 16911 1921
rect 18049 1955 18107 1961
rect 18049 1921 18061 1955
rect 18095 1921 18107 1955
rect 18049 1915 18107 1921
rect 11701 1887 11759 1893
rect 11701 1853 11713 1887
rect 11747 1853 11759 1887
rect 11701 1847 11759 1853
rect 11793 1887 11851 1893
rect 11793 1853 11805 1887
rect 11839 1884 11851 1887
rect 11974 1884 11980 1896
rect 11839 1856 11980 1884
rect 11839 1853 11851 1856
rect 11793 1847 11851 1853
rect 9398 1816 9404 1828
rect 6840 1788 9404 1816
rect 9398 1776 9404 1788
rect 9456 1776 9462 1828
rect 10318 1776 10324 1828
rect 10376 1816 10382 1828
rect 11808 1816 11836 1847
rect 11974 1844 11980 1856
rect 12032 1844 12038 1896
rect 13357 1887 13415 1893
rect 13357 1853 13369 1887
rect 13403 1884 13415 1887
rect 13403 1856 14136 1884
rect 13403 1853 13415 1856
rect 13357 1847 13415 1853
rect 13372 1816 13400 1847
rect 10376 1788 11836 1816
rect 11900 1788 13400 1816
rect 10376 1776 10382 1788
rect 6086 1708 6092 1760
rect 6144 1708 6150 1760
rect 11698 1708 11704 1760
rect 11756 1748 11762 1760
rect 11900 1748 11928 1788
rect 11756 1720 11928 1748
rect 11756 1708 11762 1720
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 14001 1751 14059 1757
rect 14001 1748 14013 1751
rect 12032 1720 14013 1748
rect 12032 1708 12038 1720
rect 14001 1717 14013 1720
rect 14047 1717 14059 1751
rect 14108 1748 14136 1856
rect 14458 1844 14464 1896
rect 14516 1884 14522 1896
rect 14737 1887 14795 1893
rect 14737 1884 14749 1887
rect 14516 1856 14749 1884
rect 14516 1844 14522 1856
rect 14737 1853 14749 1856
rect 14783 1853 14795 1887
rect 14737 1847 14795 1853
rect 15010 1844 15016 1896
rect 15068 1884 15074 1896
rect 15068 1856 15194 1884
rect 15068 1844 15074 1856
rect 15166 1816 15194 1856
rect 15838 1844 15844 1896
rect 15896 1844 15902 1896
rect 17954 1884 17960 1896
rect 17926 1844 17960 1884
rect 18012 1844 18018 1896
rect 18874 1844 18880 1896
rect 18932 1844 18938 1896
rect 17926 1816 17954 1844
rect 15166 1788 17954 1816
rect 18506 1748 18512 1760
rect 14108 1720 18512 1748
rect 14001 1711 14059 1717
rect 18506 1708 18512 1720
rect 18564 1708 18570 1760
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 5810 1504 5816 1556
rect 5868 1504 5874 1556
rect 6914 1544 6920 1556
rect 6380 1516 6920 1544
rect 5828 1476 5856 1504
rect 5460 1448 5856 1476
rect 5460 1417 5488 1448
rect 5445 1411 5503 1417
rect 5445 1377 5457 1411
rect 5491 1377 5503 1411
rect 5445 1371 5503 1377
rect 5629 1411 5687 1417
rect 5629 1377 5641 1411
rect 5675 1408 5687 1411
rect 6086 1408 6092 1420
rect 5675 1380 6092 1408
rect 5675 1377 5687 1380
rect 5629 1371 5687 1377
rect 6086 1368 6092 1380
rect 6144 1408 6150 1420
rect 6380 1417 6408 1516
rect 6914 1504 6920 1516
rect 6972 1504 6978 1556
rect 7466 1504 7472 1556
rect 7524 1504 7530 1556
rect 7926 1504 7932 1556
rect 7984 1504 7990 1556
rect 10410 1504 10416 1556
rect 10468 1544 10474 1556
rect 10965 1547 11023 1553
rect 10965 1544 10977 1547
rect 10468 1516 10977 1544
rect 10468 1504 10474 1516
rect 10965 1513 10977 1516
rect 11011 1513 11023 1547
rect 10965 1507 11023 1513
rect 7098 1476 7104 1488
rect 6656 1448 7104 1476
rect 6656 1417 6684 1448
rect 7098 1436 7104 1448
rect 7156 1436 7162 1488
rect 6181 1411 6239 1417
rect 6181 1408 6193 1411
rect 6144 1380 6193 1408
rect 6144 1368 6150 1380
rect 6181 1377 6193 1380
rect 6227 1377 6239 1411
rect 6181 1371 6239 1377
rect 6365 1411 6423 1417
rect 6365 1377 6377 1411
rect 6411 1377 6423 1411
rect 6365 1371 6423 1377
rect 6457 1411 6515 1417
rect 6457 1377 6469 1411
rect 6503 1377 6515 1411
rect 6457 1371 6515 1377
rect 6641 1411 6699 1417
rect 6641 1377 6653 1411
rect 6687 1377 6699 1411
rect 6641 1371 6699 1377
rect 6733 1411 6791 1417
rect 6733 1377 6745 1411
rect 6779 1377 6791 1411
rect 6733 1371 6791 1377
rect 6196 1340 6224 1371
rect 6472 1340 6500 1371
rect 6748 1340 6776 1371
rect 6914 1368 6920 1420
rect 6972 1368 6978 1420
rect 7009 1411 7067 1417
rect 7009 1377 7021 1411
rect 7055 1377 7067 1411
rect 7009 1371 7067 1377
rect 7024 1340 7052 1371
rect 7190 1368 7196 1420
rect 7248 1368 7254 1420
rect 7282 1368 7288 1420
rect 7340 1368 7346 1420
rect 7484 1417 7512 1504
rect 7944 1476 7972 1504
rect 11974 1476 11980 1488
rect 7944 1448 11744 1476
rect 7469 1411 7527 1417
rect 7469 1377 7481 1411
rect 7515 1377 7527 1411
rect 7469 1371 7527 1377
rect 8662 1368 8668 1420
rect 8720 1368 8726 1420
rect 9674 1368 9680 1420
rect 9732 1368 9738 1420
rect 10781 1411 10839 1417
rect 10781 1377 10793 1411
rect 10827 1377 10839 1411
rect 10781 1371 10839 1377
rect 6196 1312 7052 1340
rect 7024 1272 7052 1312
rect 7098 1300 7104 1352
rect 7156 1340 7162 1352
rect 7561 1343 7619 1349
rect 7561 1340 7573 1343
rect 7156 1312 7573 1340
rect 7156 1300 7162 1312
rect 7561 1309 7573 1312
rect 7607 1340 7619 1343
rect 7834 1340 7840 1352
rect 7607 1312 7840 1340
rect 7607 1309 7619 1312
rect 7561 1303 7619 1309
rect 7834 1300 7840 1312
rect 7892 1300 7898 1352
rect 9217 1343 9275 1349
rect 9217 1309 9229 1343
rect 9263 1340 9275 1343
rect 9692 1340 9720 1368
rect 9263 1312 9720 1340
rect 9263 1309 9275 1312
rect 9217 1303 9275 1309
rect 10686 1300 10692 1352
rect 10744 1340 10750 1352
rect 10796 1340 10824 1371
rect 11514 1368 11520 1420
rect 11572 1368 11578 1420
rect 11716 1417 11744 1448
rect 11900 1448 11980 1476
rect 11900 1417 11928 1448
rect 11974 1436 11980 1448
rect 12032 1436 12038 1488
rect 15746 1436 15752 1488
rect 15804 1436 15810 1488
rect 18506 1436 18512 1488
rect 18564 1436 18570 1488
rect 11701 1411 11759 1417
rect 11701 1377 11713 1411
rect 11747 1377 11759 1411
rect 11701 1371 11759 1377
rect 11885 1411 11943 1417
rect 11885 1377 11897 1411
rect 11931 1377 11943 1411
rect 11885 1371 11943 1377
rect 13630 1368 13636 1420
rect 13688 1408 13694 1420
rect 14829 1411 14887 1417
rect 14829 1408 14841 1411
rect 13688 1380 14841 1408
rect 13688 1368 13694 1380
rect 10744 1312 10824 1340
rect 10744 1300 10750 1312
rect 10870 1300 10876 1352
rect 10928 1340 10934 1352
rect 12069 1343 12127 1349
rect 12069 1340 12081 1343
rect 10928 1312 12081 1340
rect 10928 1300 10934 1312
rect 12069 1309 12081 1312
rect 12115 1340 12127 1343
rect 12618 1340 12624 1352
rect 12115 1312 12624 1340
rect 12115 1309 12127 1312
rect 12069 1303 12127 1309
rect 12618 1300 12624 1312
rect 12676 1340 12682 1352
rect 13446 1340 13452 1352
rect 12676 1312 13452 1340
rect 12676 1300 12682 1312
rect 13446 1300 13452 1312
rect 13504 1340 13510 1352
rect 13725 1343 13783 1349
rect 13725 1340 13737 1343
rect 13504 1312 13737 1340
rect 13504 1300 13510 1312
rect 13725 1309 13737 1312
rect 13771 1309 13783 1343
rect 13725 1303 13783 1309
rect 7282 1272 7288 1284
rect 7024 1244 7288 1272
rect 7282 1232 7288 1244
rect 7340 1232 7346 1284
rect 9030 1232 9036 1284
rect 9088 1272 9094 1284
rect 10704 1272 10732 1300
rect 9088 1244 10732 1272
rect 13541 1275 13599 1281
rect 9088 1232 9094 1244
rect 13541 1241 13553 1275
rect 13587 1272 13599 1275
rect 13832 1272 13860 1380
rect 14752 1349 14780 1380
rect 14829 1377 14841 1380
rect 14875 1377 14887 1411
rect 14829 1371 14887 1377
rect 15470 1368 15476 1420
rect 15528 1368 15534 1420
rect 17494 1368 17500 1420
rect 17552 1368 17558 1420
rect 18230 1368 18236 1420
rect 18288 1368 18294 1420
rect 19061 1411 19119 1417
rect 19061 1377 19073 1411
rect 19107 1408 19119 1411
rect 19610 1408 19616 1420
rect 19107 1380 19616 1408
rect 19107 1377 19119 1380
rect 19061 1371 19119 1377
rect 19610 1368 19616 1380
rect 19668 1368 19674 1420
rect 14737 1343 14795 1349
rect 14737 1309 14749 1343
rect 14783 1340 14795 1343
rect 14783 1312 14817 1340
rect 14783 1309 14795 1312
rect 14737 1303 14795 1309
rect 16114 1300 16120 1352
rect 16172 1340 16178 1352
rect 16393 1343 16451 1349
rect 16393 1340 16405 1343
rect 16172 1312 16405 1340
rect 16172 1300 16178 1312
rect 16393 1309 16405 1312
rect 16439 1309 16451 1343
rect 16393 1303 16451 1309
rect 17862 1300 17868 1352
rect 17920 1300 17926 1352
rect 13587 1244 13860 1272
rect 13587 1241 13599 1244
rect 13541 1235 13599 1241
rect 6086 1164 6092 1216
rect 6144 1164 6150 1216
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 6086 960 6092 1012
rect 6144 960 6150 1012
rect 6914 960 6920 1012
rect 6972 960 6978 1012
rect 7190 960 7196 1012
rect 7248 1000 7254 1012
rect 8389 1003 8447 1009
rect 8389 1000 8401 1003
rect 7248 972 8401 1000
rect 7248 960 7254 972
rect 8389 969 8401 972
rect 8435 969 8447 1003
rect 8389 963 8447 969
rect 19058 960 19064 1012
rect 19116 960 19122 1012
rect 3970 756 3976 808
rect 4028 756 4034 808
rect 5718 756 5724 808
rect 5776 796 5782 808
rect 6104 805 6132 960
rect 6932 932 6960 960
rect 8665 935 8723 941
rect 8665 932 8677 935
rect 6932 904 8677 932
rect 8665 901 8677 904
rect 8711 901 8723 935
rect 11885 935 11943 941
rect 11885 932 11897 935
rect 8665 895 8723 901
rect 9324 904 11897 932
rect 6641 867 6699 873
rect 6641 833 6653 867
rect 6687 864 6699 867
rect 7098 864 7104 876
rect 6687 836 7104 864
rect 6687 833 6699 836
rect 6641 827 6699 833
rect 7098 824 7104 836
rect 7156 824 7162 876
rect 7374 824 7380 876
rect 7432 864 7438 876
rect 8113 867 8171 873
rect 7432 836 7880 864
rect 7432 824 7438 836
rect 5813 799 5871 805
rect 5813 796 5825 799
rect 5776 768 5825 796
rect 5776 756 5782 768
rect 5813 765 5825 768
rect 5859 765 5871 799
rect 5813 759 5871 765
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 6089 799 6147 805
rect 6089 765 6101 799
rect 6135 765 6147 799
rect 6089 759 6147 765
rect 6273 799 6331 805
rect 6273 765 6285 799
rect 6319 796 6331 799
rect 6365 799 6423 805
rect 6365 796 6377 799
rect 6319 768 6377 796
rect 6319 765 6331 768
rect 6273 759 6331 765
rect 6365 765 6377 768
rect 6411 765 6423 799
rect 6365 759 6423 765
rect 6012 728 6040 759
rect 6380 728 6408 759
rect 6546 756 6552 808
rect 6604 756 6610 808
rect 7745 799 7803 805
rect 7745 765 7757 799
rect 7791 765 7803 799
rect 7852 796 7880 836
rect 8113 833 8125 867
rect 8159 864 8171 867
rect 9030 864 9036 876
rect 8159 836 9036 864
rect 8159 833 8171 836
rect 8113 827 8171 833
rect 9030 824 9036 836
rect 9088 864 9094 876
rect 9324 873 9352 904
rect 9309 867 9367 873
rect 9309 864 9321 867
rect 9088 836 9321 864
rect 9088 824 9094 836
rect 9232 805 9260 836
rect 9309 833 9321 836
rect 9355 833 9367 867
rect 9309 827 9367 833
rect 10781 867 10839 873
rect 10781 833 10793 867
rect 10827 864 10839 867
rect 10870 864 10876 876
rect 10827 836 10876 864
rect 10827 833 10839 836
rect 10781 827 10839 833
rect 10870 824 10876 836
rect 10928 824 10934 876
rect 8941 799 8999 805
rect 8941 796 8953 799
rect 7852 768 8953 796
rect 7745 759 7803 765
rect 8941 765 8953 768
rect 8987 765 8999 799
rect 8941 759 8999 765
rect 9125 799 9183 805
rect 9125 765 9137 799
rect 9171 765 9183 799
rect 9125 759 9183 765
rect 9217 799 9275 805
rect 9217 765 9229 799
rect 9263 796 9275 799
rect 9263 768 9297 796
rect 9263 765 9275 768
rect 9217 759 9275 765
rect 7760 728 7788 759
rect 8662 728 8668 740
rect 6012 700 7328 728
rect 7760 700 8668 728
rect 7300 672 7328 700
rect 8662 688 8668 700
rect 8720 688 8726 740
rect 9140 728 9168 759
rect 9398 756 9404 808
rect 9456 796 9462 808
rect 11808 805 11836 904
rect 11885 901 11897 904
rect 11931 901 11943 935
rect 11885 895 11943 901
rect 13630 892 13636 944
rect 13688 892 13694 944
rect 17589 935 17647 941
rect 17589 901 17601 935
rect 17635 932 17647 935
rect 17862 932 17868 944
rect 17635 904 17868 932
rect 17635 901 17647 904
rect 17589 895 17647 901
rect 17862 892 17868 904
rect 17920 892 17926 944
rect 13357 867 13415 873
rect 13357 833 13369 867
rect 13403 864 13415 867
rect 13446 864 13452 876
rect 13403 836 13452 864
rect 13403 833 13415 836
rect 13357 827 13415 833
rect 13446 824 13452 836
rect 13504 824 13510 876
rect 14918 824 14924 876
rect 14976 864 14982 876
rect 15105 867 15163 873
rect 15105 864 15117 867
rect 14976 836 15117 864
rect 14976 824 14982 836
rect 15105 833 15117 836
rect 15151 864 15163 867
rect 16114 864 16120 876
rect 15151 836 16120 864
rect 15151 833 15163 836
rect 15105 827 15163 833
rect 16114 824 16120 836
rect 16172 824 16178 876
rect 10965 799 11023 805
rect 10965 796 10977 799
rect 9456 768 10977 796
rect 9456 756 9462 768
rect 10965 765 10977 768
rect 11011 765 11023 799
rect 10965 759 11023 765
rect 11149 799 11207 805
rect 11149 765 11161 799
rect 11195 765 11207 799
rect 11149 759 11207 765
rect 11793 799 11851 805
rect 11793 765 11805 799
rect 11839 765 11851 799
rect 11793 759 11851 765
rect 11164 728 11192 759
rect 11974 756 11980 808
rect 12032 756 12038 808
rect 14001 799 14059 805
rect 14001 765 14013 799
rect 14047 796 14059 799
rect 15010 796 15016 808
rect 14047 768 15016 796
rect 14047 765 14059 768
rect 14001 759 14059 765
rect 15010 756 15016 768
rect 15068 756 15074 808
rect 17494 756 17500 808
rect 17552 756 17558 808
rect 11992 728 12020 756
rect 9140 700 12020 728
rect 7282 620 7288 672
rect 7340 660 7346 672
rect 9140 660 9168 700
rect 7340 632 9168 660
rect 7340 620 7346 632
rect 15470 620 15476 672
rect 15528 660 15534 672
rect 17773 663 17831 669
rect 17773 660 17785 663
rect 15528 632 17785 660
rect 15528 620 15534 632
rect 17773 629 17785 632
rect 17819 629 17831 663
rect 17773 623 17831 629
rect 18046 620 18052 672
rect 18104 660 18110 672
rect 18325 663 18383 669
rect 18325 660 18337 663
rect 18104 632 18337 660
rect 18104 620 18110 632
rect 18325 629 18337 632
rect 18371 629 18383 663
rect 18325 623 18383 629
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 3884 18912 3936 18964
rect 7748 18844 7800 18896
rect 8116 18776 8168 18828
rect 15476 18776 15528 18828
rect 16120 18776 16172 18828
rect 18052 18776 18104 18828
rect 848 18751 900 18760
rect 848 18717 857 18751
rect 857 18717 891 18751
rect 891 18717 900 18751
rect 848 18708 900 18717
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 9680 18708 9732 18760
rect 10416 18708 10468 18760
rect 8668 18683 8720 18692
rect 8668 18649 8677 18683
rect 8677 18649 8711 18683
rect 8711 18649 8720 18683
rect 8668 18640 8720 18649
rect 9680 18572 9732 18624
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 10508 18232 10560 18284
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 6092 18096 6144 18148
rect 8944 18096 8996 18148
rect 10232 18096 10284 18148
rect 6828 18028 6880 18080
rect 8116 18071 8168 18080
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 9220 18028 9272 18080
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 4896 17756 4948 17808
rect 7288 17824 7340 17876
rect 9680 17824 9732 17876
rect 10232 17824 10284 17876
rect 5448 17688 5500 17740
rect 5724 17688 5776 17740
rect 7104 17756 7156 17808
rect 7380 17756 7432 17808
rect 8944 17688 8996 17740
rect 12532 17756 12584 17808
rect 10968 17731 11020 17740
rect 10968 17697 10977 17731
rect 10977 17697 11011 17731
rect 11011 17697 11020 17731
rect 10968 17688 11020 17697
rect 3516 17620 3568 17672
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 6368 17620 6420 17672
rect 8852 17620 8904 17672
rect 10508 17620 10560 17672
rect 5816 17527 5868 17536
rect 5816 17493 5825 17527
rect 5825 17493 5859 17527
rect 5859 17493 5868 17527
rect 5816 17484 5868 17493
rect 6368 17484 6420 17536
rect 6828 17484 6880 17536
rect 7196 17484 7248 17536
rect 11888 17484 11940 17536
rect 12624 17484 12676 17536
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 3884 17280 3936 17332
rect 5816 17280 5868 17332
rect 6092 17323 6144 17332
rect 6092 17289 6101 17323
rect 6101 17289 6135 17323
rect 6135 17289 6144 17323
rect 6092 17280 6144 17289
rect 5448 17212 5500 17264
rect 6368 17212 6420 17264
rect 7380 17280 7432 17332
rect 10968 17280 11020 17332
rect 5448 17076 5500 17128
rect 6276 17119 6328 17128
rect 6276 17085 6285 17119
rect 6285 17085 6319 17119
rect 6319 17085 6328 17119
rect 6276 17076 6328 17085
rect 5540 17008 5592 17060
rect 5632 17008 5684 17060
rect 6644 17119 6696 17128
rect 6644 17085 6653 17119
rect 6653 17085 6687 17119
rect 6687 17085 6696 17119
rect 6644 17076 6696 17085
rect 7104 17144 7156 17196
rect 7288 17076 7340 17128
rect 5724 16940 5776 16992
rect 7104 16940 7156 16992
rect 7196 16940 7248 16992
rect 7380 16940 7432 16992
rect 8760 17119 8812 17128
rect 8760 17085 8769 17119
rect 8769 17085 8803 17119
rect 8803 17085 8812 17119
rect 8760 17076 8812 17085
rect 8852 17076 8904 17128
rect 10508 17144 10560 17196
rect 11704 17144 11756 17196
rect 12624 17076 12676 17128
rect 7564 17008 7616 17060
rect 12532 17008 12584 17060
rect 9680 16940 9732 16992
rect 10600 16940 10652 16992
rect 11888 16940 11940 16992
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 6644 16736 6696 16788
rect 3700 16643 3752 16652
rect 3700 16609 3709 16643
rect 3709 16609 3743 16643
rect 3743 16609 3752 16643
rect 3700 16600 3752 16609
rect 5540 16600 5592 16652
rect 6184 16600 6236 16652
rect 6920 16668 6972 16720
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 7104 16779 7156 16788
rect 7104 16745 7113 16779
rect 7113 16745 7147 16779
rect 7147 16745 7156 16779
rect 7104 16736 7156 16745
rect 8760 16736 8812 16788
rect 9680 16736 9732 16788
rect 7196 16668 7248 16720
rect 7380 16668 7432 16720
rect 5908 16532 5960 16584
rect 15752 16600 15804 16652
rect 18972 16643 19024 16652
rect 18972 16609 18981 16643
rect 18981 16609 19015 16643
rect 19015 16609 19024 16643
rect 18972 16600 19024 16609
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 3424 16396 3476 16448
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 6828 16396 6880 16448
rect 7564 16396 7616 16448
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 3976 16192 4028 16244
rect 6644 16192 6696 16244
rect 6920 16192 6972 16244
rect 4988 16167 5040 16176
rect 4988 16133 4997 16167
rect 4997 16133 5031 16167
rect 5031 16133 5040 16167
rect 4988 16124 5040 16133
rect 3516 16056 3568 16108
rect 8852 16056 8904 16108
rect 9128 16056 9180 16108
rect 11428 16056 11480 16108
rect 3424 15920 3476 15972
rect 4344 15852 4396 15904
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 11704 16056 11756 16108
rect 12072 15988 12124 16040
rect 19064 15988 19116 16040
rect 5724 15852 5776 15904
rect 7840 15852 7892 15904
rect 8300 15852 8352 15904
rect 8484 15852 8536 15904
rect 9220 15852 9272 15904
rect 10692 15920 10744 15972
rect 11520 15920 11572 15972
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 11612 15852 11664 15861
rect 12256 15852 12308 15904
rect 16580 15852 16632 15904
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 3884 15580 3936 15632
rect 3976 15623 4028 15632
rect 3976 15589 3985 15623
rect 3985 15589 4019 15623
rect 4019 15589 4028 15623
rect 3976 15580 4028 15589
rect 3148 15512 3200 15564
rect 3700 15444 3752 15496
rect 5448 15648 5500 15700
rect 5724 15580 5776 15632
rect 5632 15512 5684 15564
rect 5908 15691 5960 15700
rect 5908 15657 5917 15691
rect 5917 15657 5951 15691
rect 5951 15657 5960 15691
rect 5908 15648 5960 15657
rect 6368 15623 6420 15632
rect 6368 15589 6377 15623
rect 6377 15589 6411 15623
rect 6411 15589 6420 15623
rect 6368 15580 6420 15589
rect 9128 15648 9180 15700
rect 8208 15623 8260 15632
rect 8208 15589 8217 15623
rect 8217 15589 8251 15623
rect 8251 15589 8260 15623
rect 8208 15580 8260 15589
rect 8944 15580 8996 15632
rect 9588 15648 9640 15700
rect 11244 15648 11296 15700
rect 11612 15648 11664 15700
rect 11704 15648 11756 15700
rect 12072 15648 12124 15700
rect 6000 15555 6052 15564
rect 6000 15521 6009 15555
rect 6009 15521 6043 15555
rect 6043 15521 6052 15555
rect 6000 15512 6052 15521
rect 6092 15555 6144 15564
rect 6092 15521 6101 15555
rect 6101 15521 6135 15555
rect 6135 15521 6144 15555
rect 6092 15512 6144 15521
rect 4620 15444 4672 15496
rect 4068 15376 4120 15428
rect 5908 15444 5960 15496
rect 6736 15444 6788 15496
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 9588 15512 9640 15564
rect 10232 15512 10284 15564
rect 8944 15444 8996 15496
rect 9220 15444 9272 15496
rect 1860 15308 1912 15360
rect 5172 15308 5224 15360
rect 6552 15308 6604 15360
rect 7840 15351 7892 15360
rect 7840 15317 7849 15351
rect 7849 15317 7883 15351
rect 7883 15317 7892 15351
rect 12256 15580 12308 15632
rect 12532 15580 12584 15632
rect 11428 15512 11480 15564
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 18328 15444 18380 15496
rect 7840 15308 7892 15317
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 3516 15104 3568 15156
rect 3884 15147 3936 15156
rect 3884 15113 3893 15147
rect 3893 15113 3927 15147
rect 3927 15113 3936 15147
rect 3884 15104 3936 15113
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 4896 15104 4948 15156
rect 4804 15036 4856 15088
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 3148 14968 3200 15020
rect 3976 14968 4028 15020
rect 848 14943 900 14952
rect 848 14909 857 14943
rect 857 14909 891 14943
rect 891 14909 900 14943
rect 848 14900 900 14909
rect 1124 14875 1176 14884
rect 1124 14841 1133 14875
rect 1133 14841 1167 14875
rect 1167 14841 1176 14875
rect 1124 14832 1176 14841
rect 2688 14832 2740 14884
rect 3424 14900 3476 14952
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4896 14900 4948 14952
rect 6736 15104 6788 15156
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 8208 15147 8260 15156
rect 8208 15113 8217 15147
rect 8217 15113 8251 15147
rect 8251 15113 8260 15147
rect 8208 15104 8260 15113
rect 8484 15036 8536 15088
rect 8944 15036 8996 15088
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 18328 15079 18380 15088
rect 18328 15045 18337 15079
rect 18337 15045 18371 15079
rect 18371 15045 18380 15079
rect 18328 15036 18380 15045
rect 6920 14900 6972 14952
rect 4988 14832 5040 14884
rect 5172 14832 5224 14884
rect 8300 14900 8352 14952
rect 8944 14900 8996 14952
rect 12532 14968 12584 15020
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 11428 14900 11480 14952
rect 16948 14968 17000 15020
rect 17500 14968 17552 15020
rect 7288 14832 7340 14884
rect 3148 14764 3200 14816
rect 7104 14764 7156 14816
rect 9404 14875 9456 14884
rect 9404 14841 9413 14875
rect 9413 14841 9447 14875
rect 9447 14841 9456 14875
rect 9404 14832 9456 14841
rect 10692 14764 10744 14816
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 15844 14832 15896 14884
rect 19064 14832 19116 14884
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 1124 14560 1176 14612
rect 2412 14560 2464 14612
rect 3516 14560 3568 14612
rect 4068 14560 4120 14612
rect 4896 14560 4948 14612
rect 5448 14560 5500 14612
rect 7012 14560 7064 14612
rect 7932 14560 7984 14612
rect 8944 14560 8996 14612
rect 9404 14560 9456 14612
rect 11336 14560 11388 14612
rect 14924 14603 14976 14612
rect 14924 14569 14933 14603
rect 14933 14569 14967 14603
rect 14967 14569 14976 14603
rect 14924 14560 14976 14569
rect 2872 14492 2924 14544
rect 4160 14492 4212 14544
rect 5632 14492 5684 14544
rect 6000 14492 6052 14544
rect 6736 14492 6788 14544
rect 15016 14535 15068 14544
rect 15016 14501 15025 14535
rect 15025 14501 15059 14535
rect 15059 14501 15068 14535
rect 15016 14492 15068 14501
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 2044 14424 2096 14476
rect 2320 14467 2372 14476
rect 2320 14433 2329 14467
rect 2329 14433 2363 14467
rect 2363 14433 2372 14467
rect 2320 14424 2372 14433
rect 2136 14356 2188 14408
rect 848 14220 900 14272
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 2688 14356 2740 14408
rect 4344 14424 4396 14476
rect 4988 14424 5040 14476
rect 5448 14424 5500 14476
rect 7012 14424 7064 14476
rect 9680 14424 9732 14476
rect 11980 14424 12032 14476
rect 13084 14424 13136 14476
rect 13360 14424 13412 14476
rect 4252 14331 4304 14340
rect 4252 14297 4261 14331
rect 4261 14297 4295 14331
rect 4295 14297 4304 14331
rect 4252 14288 4304 14297
rect 11704 14356 11756 14408
rect 12532 14356 12584 14408
rect 15292 14424 15344 14476
rect 15844 14424 15896 14476
rect 16580 14492 16632 14544
rect 15200 14356 15252 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 6184 14288 6236 14340
rect 10140 14288 10192 14340
rect 10692 14288 10744 14340
rect 10876 14288 10928 14340
rect 5908 14220 5960 14272
rect 10600 14220 10652 14272
rect 12900 14288 12952 14340
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 17316 14424 17368 14476
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 18880 14356 18932 14408
rect 17592 14288 17644 14340
rect 18328 14288 18380 14340
rect 12992 14220 13044 14272
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 18696 14263 18748 14272
rect 18696 14229 18705 14263
rect 18705 14229 18739 14263
rect 18739 14229 18748 14263
rect 18696 14220 18748 14229
rect 18972 14220 19024 14272
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 2136 14016 2188 14068
rect 2596 14016 2648 14068
rect 4804 14016 4856 14068
rect 6000 14016 6052 14068
rect 9680 14016 9732 14068
rect 9772 14016 9824 14068
rect 7380 13948 7432 14000
rect 7840 13948 7892 14000
rect 3148 13880 3200 13932
rect 2044 13744 2096 13796
rect 5540 13880 5592 13932
rect 6644 13880 6696 13932
rect 10140 13880 10192 13932
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 4252 13812 4304 13864
rect 7012 13812 7064 13864
rect 7104 13812 7156 13864
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 7472 13812 7524 13864
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 10232 13855 10284 13864
rect 10232 13821 10241 13855
rect 10241 13821 10275 13855
rect 10275 13821 10284 13855
rect 10232 13812 10284 13821
rect 10968 14016 11020 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 11060 13948 11112 14000
rect 15016 13948 15068 14000
rect 15292 13948 15344 14000
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 6552 13787 6604 13796
rect 6552 13753 6561 13787
rect 6561 13753 6595 13787
rect 6595 13753 6604 13787
rect 6552 13744 6604 13753
rect 9128 13744 9180 13796
rect 6828 13676 6880 13728
rect 7104 13676 7156 13728
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 12624 13812 12676 13864
rect 14464 13812 14516 13864
rect 14924 13812 14976 13864
rect 16212 13812 16264 13864
rect 17592 13812 17644 13864
rect 18880 13812 18932 13864
rect 19156 13812 19208 13864
rect 11428 13744 11480 13796
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 11336 13676 11388 13728
rect 12348 13744 12400 13796
rect 13360 13744 13412 13796
rect 15200 13744 15252 13796
rect 15568 13744 15620 13796
rect 12808 13676 12860 13728
rect 18696 13676 18748 13728
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 4988 13472 5040 13524
rect 6000 13515 6052 13524
rect 6000 13481 6027 13515
rect 6027 13481 6052 13515
rect 6000 13472 6052 13481
rect 4252 13404 4304 13456
rect 5356 13404 5408 13456
rect 7472 13472 7524 13524
rect 2136 13336 2188 13388
rect 3148 13336 3200 13388
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2044 13268 2096 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 6736 13404 6788 13456
rect 7104 13404 7156 13456
rect 7288 13404 7340 13456
rect 6092 13336 6144 13388
rect 4896 13268 4948 13277
rect 6828 13268 6880 13320
rect 8300 13336 8352 13388
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 9128 13447 9180 13456
rect 9128 13413 9137 13447
rect 9137 13413 9171 13447
rect 9171 13413 9180 13447
rect 9128 13404 9180 13413
rect 8208 13268 8260 13320
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 4528 13200 4580 13252
rect 1768 13175 1820 13184
rect 1768 13141 1777 13175
rect 1777 13141 1811 13175
rect 1811 13141 1820 13175
rect 1768 13132 1820 13141
rect 3516 13132 3568 13184
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 5448 13132 5500 13141
rect 8116 13132 8168 13184
rect 8944 13200 8996 13252
rect 9496 13336 9548 13388
rect 10692 13404 10744 13456
rect 12348 13472 12400 13524
rect 14096 13472 14148 13524
rect 10876 13336 10928 13388
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 11244 13379 11296 13388
rect 11244 13345 11254 13379
rect 11254 13345 11288 13379
rect 11288 13345 11296 13379
rect 11244 13336 11296 13345
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 10232 13268 10284 13320
rect 10508 13268 10560 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11520 13379 11572 13388
rect 11520 13345 11529 13379
rect 11529 13345 11563 13379
rect 11563 13345 11572 13379
rect 11520 13336 11572 13345
rect 11704 13336 11756 13388
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 12532 13336 12584 13388
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 13176 13379 13228 13388
rect 13176 13345 13211 13379
rect 13211 13345 13228 13379
rect 13176 13336 13228 13345
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 14464 13379 14516 13388
rect 14464 13345 14473 13379
rect 14473 13345 14507 13379
rect 14507 13345 14516 13379
rect 14464 13336 14516 13345
rect 9864 13200 9916 13252
rect 14280 13243 14332 13252
rect 14280 13209 14289 13243
rect 14289 13209 14323 13243
rect 14323 13209 14332 13243
rect 17500 13472 17552 13524
rect 15016 13379 15068 13388
rect 15016 13345 15025 13379
rect 15025 13345 15059 13379
rect 15059 13345 15068 13379
rect 15016 13336 15068 13345
rect 15292 13336 15344 13388
rect 15568 13379 15620 13388
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 15568 13336 15620 13345
rect 16212 13404 16264 13456
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 18236 13379 18288 13388
rect 18236 13345 18245 13379
rect 18245 13345 18279 13379
rect 18279 13345 18288 13379
rect 18236 13336 18288 13345
rect 14280 13200 14332 13209
rect 17868 13200 17920 13252
rect 9312 13132 9364 13184
rect 10968 13132 11020 13184
rect 11980 13132 12032 13184
rect 12532 13132 12584 13184
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13820 13132 13872 13184
rect 14556 13175 14608 13184
rect 14556 13141 14565 13175
rect 14565 13141 14599 13175
rect 14599 13141 14608 13175
rect 14556 13132 14608 13141
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 3148 12860 3200 12912
rect 1768 12792 1820 12844
rect 848 12767 900 12776
rect 848 12733 857 12767
rect 857 12733 891 12767
rect 891 12733 900 12767
rect 848 12724 900 12733
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 3700 12767 3752 12776
rect 3700 12733 3709 12767
rect 3709 12733 3743 12767
rect 3743 12733 3752 12767
rect 3700 12724 3752 12733
rect 3976 12724 4028 12776
rect 2504 12656 2556 12708
rect 2688 12699 2740 12708
rect 2688 12665 2697 12699
rect 2697 12665 2731 12699
rect 2731 12665 2740 12699
rect 2688 12656 2740 12665
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 3792 12588 3844 12640
rect 4160 12792 4212 12844
rect 4804 12928 4856 12980
rect 5172 12928 5224 12980
rect 7196 12971 7248 12980
rect 7196 12937 7205 12971
rect 7205 12937 7239 12971
rect 7239 12937 7248 12971
rect 7196 12928 7248 12937
rect 8668 12928 8720 12980
rect 4988 12792 5040 12844
rect 5264 12792 5316 12844
rect 4344 12656 4396 12708
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 8116 12860 8168 12912
rect 9404 12860 9456 12912
rect 9496 12860 9548 12912
rect 6828 12792 6880 12801
rect 7196 12724 7248 12776
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 8484 12724 8536 12776
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 8852 12792 8904 12844
rect 8944 12792 8996 12844
rect 10324 12928 10376 12980
rect 9772 12792 9824 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 9220 12724 9272 12776
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 9404 12724 9456 12776
rect 11336 12928 11388 12980
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 12532 12971 12584 12980
rect 12532 12937 12541 12971
rect 12541 12937 12575 12971
rect 12575 12937 12584 12971
rect 12532 12928 12584 12937
rect 12716 12928 12768 12980
rect 10692 12860 10744 12912
rect 10876 12860 10928 12912
rect 10784 12792 10836 12844
rect 12348 12860 12400 12912
rect 12992 12860 13044 12912
rect 13820 12860 13872 12912
rect 14096 12835 14148 12844
rect 14096 12801 14114 12835
rect 14114 12801 14148 12835
rect 14096 12792 14148 12801
rect 14280 12792 14332 12844
rect 15568 12860 15620 12912
rect 16212 12835 16264 12844
rect 16212 12801 16221 12835
rect 16221 12801 16255 12835
rect 16255 12801 16264 12835
rect 16212 12792 16264 12801
rect 11060 12724 11112 12776
rect 11520 12724 11572 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 16488 12724 16540 12776
rect 18604 12792 18656 12844
rect 5264 12588 5316 12640
rect 5356 12588 5408 12640
rect 7840 12588 7892 12640
rect 10784 12699 10836 12708
rect 10784 12665 10793 12699
rect 10793 12665 10827 12699
rect 10827 12665 10836 12699
rect 10784 12656 10836 12665
rect 9128 12588 9180 12640
rect 9496 12588 9548 12640
rect 9588 12588 9640 12640
rect 9772 12588 9824 12640
rect 10508 12588 10560 12640
rect 12072 12588 12124 12640
rect 12532 12588 12584 12640
rect 13544 12699 13596 12708
rect 13544 12665 13553 12699
rect 13553 12665 13587 12699
rect 13587 12665 13596 12699
rect 13544 12656 13596 12665
rect 15292 12588 15344 12640
rect 17868 12588 17920 12640
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 1676 12248 1728 12300
rect 2688 12359 2740 12368
rect 2688 12325 2697 12359
rect 2697 12325 2731 12359
rect 2731 12325 2740 12359
rect 2688 12316 2740 12325
rect 2136 12180 2188 12232
rect 1860 12112 1912 12164
rect 2412 12180 2464 12232
rect 3700 12384 3752 12436
rect 3792 12384 3844 12436
rect 4896 12427 4948 12436
rect 4896 12393 4905 12427
rect 4905 12393 4939 12427
rect 4939 12393 4948 12427
rect 4896 12384 4948 12393
rect 8208 12384 8260 12436
rect 3424 12359 3476 12368
rect 3424 12325 3433 12359
rect 3433 12325 3467 12359
rect 3467 12325 3476 12359
rect 3424 12316 3476 12325
rect 4436 12248 4488 12300
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 6644 12248 6696 12300
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 10600 12384 10652 12436
rect 11612 12384 11664 12436
rect 12624 12384 12676 12436
rect 12900 12384 12952 12436
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 9036 12359 9088 12368
rect 9036 12325 9045 12359
rect 9045 12325 9079 12359
rect 9079 12325 9088 12359
rect 9036 12316 9088 12325
rect 9128 12316 9180 12368
rect 11060 12316 11112 12368
rect 11244 12316 11296 12368
rect 12164 12359 12216 12368
rect 12164 12325 12173 12359
rect 12173 12325 12207 12359
rect 12207 12325 12216 12359
rect 12164 12316 12216 12325
rect 15200 12384 15252 12436
rect 16672 12384 16724 12436
rect 9220 12248 9272 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 11428 12291 11480 12300
rect 11428 12257 11437 12291
rect 11437 12257 11471 12291
rect 11471 12257 11480 12291
rect 11428 12248 11480 12257
rect 11796 12248 11848 12300
rect 3056 12112 3108 12164
rect 2596 12044 2648 12096
rect 9128 12112 9180 12164
rect 9312 12112 9364 12164
rect 9680 12112 9732 12164
rect 11060 12112 11112 12164
rect 4160 12044 4212 12096
rect 6184 12044 6236 12096
rect 9220 12044 9272 12096
rect 10324 12044 10376 12096
rect 10784 12044 10836 12096
rect 12348 12248 12400 12300
rect 12256 12155 12308 12164
rect 12256 12121 12265 12155
rect 12265 12121 12299 12155
rect 12299 12121 12308 12155
rect 12256 12112 12308 12121
rect 13820 12316 13872 12368
rect 15108 12248 15160 12300
rect 15568 12248 15620 12300
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 13360 12223 13412 12232
rect 13360 12189 13378 12223
rect 13378 12189 13412 12223
rect 13360 12180 13412 12189
rect 14004 12180 14056 12232
rect 15292 12180 15344 12232
rect 12716 12044 12768 12096
rect 15108 12112 15160 12164
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 18880 12180 18932 12232
rect 17868 12112 17920 12164
rect 13360 12044 13412 12096
rect 16304 12044 16356 12096
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 1492 11815 1544 11824
rect 1492 11781 1501 11815
rect 1501 11781 1535 11815
rect 1535 11781 1544 11815
rect 1492 11772 1544 11781
rect 3332 11772 3384 11824
rect 1584 11636 1636 11688
rect 2412 11636 2464 11688
rect 3240 11636 3292 11688
rect 4804 11840 4856 11892
rect 7564 11883 7616 11892
rect 7564 11849 7573 11883
rect 7573 11849 7607 11883
rect 7607 11849 7616 11883
rect 7564 11840 7616 11849
rect 10416 11840 10468 11892
rect 12440 11772 12492 11824
rect 13084 11772 13136 11824
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6184 11704 6236 11756
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 10048 11704 10100 11756
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 4988 11636 5040 11688
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 11060 11679 11112 11688
rect 1676 11500 1728 11552
rect 2596 11500 2648 11552
rect 4620 11568 4672 11620
rect 6552 11568 6604 11620
rect 8944 11568 8996 11620
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 11244 11679 11296 11688
rect 11244 11645 11253 11679
rect 11253 11645 11287 11679
rect 11287 11645 11296 11679
rect 11244 11636 11296 11645
rect 11428 11636 11480 11688
rect 11704 11636 11756 11688
rect 12808 11636 12860 11688
rect 13544 11636 13596 11688
rect 15108 11704 15160 11756
rect 15292 11636 15344 11688
rect 16488 11636 16540 11688
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 17868 11636 17920 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 4436 11500 4488 11552
rect 4804 11500 4856 11552
rect 5448 11500 5500 11552
rect 8116 11500 8168 11552
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 9128 11500 9180 11552
rect 9404 11500 9456 11552
rect 11520 11568 11572 11620
rect 15108 11568 15160 11620
rect 17132 11611 17184 11620
rect 17132 11577 17141 11611
rect 17141 11577 17175 11611
rect 17175 11577 17184 11611
rect 17132 11568 17184 11577
rect 10784 11500 10836 11552
rect 12624 11500 12676 11552
rect 13360 11500 13412 11552
rect 14188 11500 14240 11552
rect 15016 11500 15068 11552
rect 17316 11500 17368 11552
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 2504 11228 2556 11280
rect 848 11203 900 11212
rect 848 11169 857 11203
rect 857 11169 891 11203
rect 891 11169 900 11203
rect 848 11160 900 11169
rect 4160 11296 4212 11348
rect 4988 11296 5040 11348
rect 5448 11296 5500 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 7564 11296 7616 11348
rect 8668 11296 8720 11348
rect 8852 11296 8904 11348
rect 9036 11296 9088 11348
rect 9404 11296 9456 11348
rect 9680 11296 9732 11348
rect 4436 11228 4488 11280
rect 6552 11228 6604 11280
rect 6000 11160 6052 11212
rect 1124 11135 1176 11144
rect 1124 11101 1133 11135
rect 1133 11101 1167 11135
rect 1167 11101 1176 11135
rect 1124 11092 1176 11101
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 6828 11092 6880 11144
rect 4620 11067 4672 11076
rect 4620 11033 4629 11067
rect 4629 11033 4663 11067
rect 4663 11033 4672 11067
rect 7380 11228 7432 11280
rect 7196 11160 7248 11212
rect 8392 11228 8444 11280
rect 4620 11024 4672 11033
rect 2412 10956 2464 11008
rect 5448 10956 5500 11008
rect 8300 11160 8352 11212
rect 10232 11296 10284 11348
rect 11060 11296 11112 11348
rect 12440 11296 12492 11348
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 10692 11228 10744 11280
rect 10784 11228 10836 11280
rect 9128 11092 9180 11144
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10232 11203 10284 11212
rect 10232 11169 10249 11203
rect 10249 11169 10284 11203
rect 10232 11160 10284 11169
rect 8576 11024 8628 11076
rect 9956 11092 10008 11144
rect 11520 11160 11572 11212
rect 9588 11024 9640 11076
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 17408 11296 17460 11348
rect 13360 11271 13412 11280
rect 13360 11237 13369 11271
rect 13369 11237 13403 11271
rect 13403 11237 13412 11271
rect 13360 11228 13412 11237
rect 13820 11271 13872 11280
rect 13820 11237 13829 11271
rect 13829 11237 13863 11271
rect 13863 11237 13872 11271
rect 13820 11228 13872 11237
rect 15292 11228 15344 11280
rect 18236 11228 18288 11280
rect 18880 11271 18932 11280
rect 18880 11237 18889 11271
rect 18889 11237 18923 11271
rect 18923 11237 18932 11271
rect 18880 11228 18932 11237
rect 12808 11160 12860 11212
rect 12992 11203 13044 11212
rect 12992 11169 13001 11203
rect 13001 11169 13035 11203
rect 13035 11169 13044 11203
rect 12992 11160 13044 11169
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 15200 11160 15252 11212
rect 16488 11203 16540 11212
rect 16488 11169 16497 11203
rect 16497 11169 16531 11203
rect 16531 11169 16540 11203
rect 16488 11160 16540 11169
rect 10232 11024 10284 11076
rect 10600 11024 10652 11076
rect 10692 11067 10744 11076
rect 10692 11033 10701 11067
rect 10701 11033 10735 11067
rect 10735 11033 10744 11067
rect 10692 11024 10744 11033
rect 11612 11024 11664 11076
rect 9864 10956 9916 11008
rect 10140 10956 10192 11008
rect 10784 10956 10836 11008
rect 13820 11067 13872 11076
rect 13820 11033 13829 11067
rect 13829 11033 13863 11067
rect 13863 11033 13872 11067
rect 13820 11024 13872 11033
rect 13912 11024 13964 11076
rect 14832 11024 14884 11076
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 17868 11024 17920 11076
rect 17132 10956 17184 11008
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 1124 10752 1176 10804
rect 3148 10752 3200 10804
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 9312 10752 9364 10804
rect 9404 10752 9456 10804
rect 3332 10727 3384 10736
rect 3332 10693 3341 10727
rect 3341 10693 3375 10727
rect 3375 10693 3384 10727
rect 3332 10684 3384 10693
rect 8760 10684 8812 10736
rect 2412 10616 2464 10668
rect 1492 10591 1544 10600
rect 1492 10557 1501 10591
rect 1501 10557 1535 10591
rect 1535 10557 1544 10591
rect 1492 10548 1544 10557
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 3516 10616 3568 10668
rect 4160 10616 4212 10668
rect 5816 10616 5868 10668
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 6552 10548 6604 10600
rect 8576 10548 8628 10600
rect 8668 10548 8720 10600
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 10140 10684 10192 10736
rect 9864 10616 9916 10668
rect 10048 10616 10100 10668
rect 11612 10752 11664 10804
rect 11336 10684 11388 10736
rect 13912 10684 13964 10736
rect 14924 10684 14976 10736
rect 15016 10616 15068 10668
rect 15292 10616 15344 10668
rect 3424 10412 3476 10464
rect 4804 10480 4856 10532
rect 8760 10412 8812 10464
rect 8944 10412 8996 10464
rect 10324 10480 10376 10532
rect 10784 10548 10836 10600
rect 14004 10548 14056 10600
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 14924 10548 14976 10600
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15568 10616 15620 10668
rect 16488 10616 16540 10668
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 15200 10548 15252 10557
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 17960 10591 18012 10600
rect 17960 10557 17969 10591
rect 17969 10557 18003 10591
rect 18003 10557 18012 10591
rect 17960 10548 18012 10557
rect 18696 10548 18748 10600
rect 10876 10480 10928 10532
rect 13820 10480 13872 10532
rect 14188 10480 14240 10532
rect 9956 10412 10008 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 15108 10412 15160 10464
rect 15936 10523 15988 10532
rect 15936 10489 15945 10523
rect 15945 10489 15979 10523
rect 15979 10489 15988 10523
rect 15936 10480 15988 10489
rect 16212 10480 16264 10532
rect 16488 10412 16540 10464
rect 17408 10412 17460 10464
rect 18144 10412 18196 10464
rect 19064 10412 19116 10464
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 3148 10208 3200 10260
rect 2596 10140 2648 10192
rect 3608 10140 3660 10192
rect 7288 10140 7340 10192
rect 2504 10072 2556 10124
rect 3240 10072 3292 10124
rect 8392 10072 8444 10124
rect 9220 10072 9272 10124
rect 9956 10208 10008 10260
rect 11336 10208 11388 10260
rect 10600 10140 10652 10192
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 10232 10072 10284 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 3516 9936 3568 9988
rect 3884 9936 3936 9988
rect 6368 9868 6420 9920
rect 7012 9868 7064 9920
rect 7932 9868 7984 9920
rect 10048 10004 10100 10056
rect 10876 10072 10928 10124
rect 11244 10072 11296 10124
rect 11520 10072 11572 10124
rect 12440 10072 12492 10124
rect 13820 10208 13872 10260
rect 14188 10208 14240 10260
rect 15200 10208 15252 10260
rect 15384 10251 15436 10260
rect 15384 10217 15393 10251
rect 15393 10217 15427 10251
rect 15427 10217 15436 10251
rect 15384 10208 15436 10217
rect 15936 10208 15988 10260
rect 12808 10072 12860 10124
rect 12624 10004 12676 10056
rect 12992 10004 13044 10056
rect 10140 9936 10192 9988
rect 10232 9936 10284 9988
rect 10968 9868 11020 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11704 9868 11756 9920
rect 12440 9868 12492 9920
rect 13820 10072 13872 10124
rect 14188 10072 14240 10124
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 15200 10115 15252 10124
rect 15200 10081 15209 10115
rect 15209 10081 15243 10115
rect 15243 10081 15252 10115
rect 15200 10072 15252 10081
rect 13912 9936 13964 9988
rect 14464 10047 14516 10056
rect 14464 10013 14498 10047
rect 14498 10013 14516 10047
rect 14464 10004 14516 10013
rect 15108 10004 15160 10056
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 16488 10115 16540 10124
rect 16488 10081 16497 10115
rect 16497 10081 16531 10115
rect 16531 10081 16540 10115
rect 16488 10072 16540 10081
rect 16580 10072 16632 10124
rect 16764 10115 16816 10124
rect 16764 10081 16773 10115
rect 16773 10081 16807 10115
rect 16807 10081 16816 10115
rect 16764 10072 16816 10081
rect 17224 10072 17276 10124
rect 17500 10072 17552 10124
rect 15016 9936 15068 9988
rect 15200 9936 15252 9988
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 13268 9868 13320 9877
rect 14648 9911 14700 9920
rect 14648 9877 14657 9911
rect 14657 9877 14691 9911
rect 14691 9877 14700 9911
rect 14648 9868 14700 9877
rect 14924 9868 14976 9920
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17960 10004 18012 10056
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 15568 9936 15620 9988
rect 16120 9979 16172 9988
rect 16120 9945 16129 9979
rect 16129 9945 16163 9979
rect 16163 9945 16172 9979
rect 16120 9936 16172 9945
rect 18512 9936 18564 9988
rect 15844 9868 15896 9920
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 16396 9868 16448 9877
rect 18972 9868 19024 9920
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 9864 9664 9916 9716
rect 1676 9596 1728 9648
rect 10600 9664 10652 9716
rect 10968 9664 11020 9716
rect 10692 9596 10744 9648
rect 5816 9528 5868 9580
rect 6368 9528 6420 9580
rect 8760 9528 8812 9580
rect 1952 9460 2004 9512
rect 2504 9460 2556 9512
rect 3148 9460 3200 9512
rect 8392 9460 8444 9512
rect 9128 9528 9180 9580
rect 9312 9528 9364 9580
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 10600 9528 10652 9580
rect 10140 9460 10192 9512
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 10416 9503 10468 9512
rect 10416 9469 10423 9503
rect 10423 9469 10468 9503
rect 10416 9460 10468 9469
rect 10508 9503 10560 9512
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 10876 9460 10928 9512
rect 11152 9528 11204 9580
rect 11428 9528 11480 9580
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 6736 9392 6788 9444
rect 9680 9392 9732 9444
rect 1584 9324 1636 9376
rect 3516 9324 3568 9376
rect 4252 9324 4304 9376
rect 7288 9324 7340 9376
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 9128 9324 9180 9376
rect 11336 9503 11388 9512
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 11888 9528 11940 9580
rect 12992 9664 13044 9716
rect 14464 9664 14516 9716
rect 15660 9664 15712 9716
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 18696 9707 18748 9716
rect 18696 9673 18705 9707
rect 18705 9673 18739 9707
rect 18739 9673 18748 9707
rect 18696 9664 18748 9673
rect 14096 9596 14148 9648
rect 18052 9596 18104 9648
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 11612 9392 11664 9444
rect 12716 9528 12768 9580
rect 12808 9528 12860 9580
rect 12900 9528 12952 9580
rect 15200 9528 15252 9580
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 14372 9460 14424 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 11796 9324 11848 9376
rect 12532 9324 12584 9376
rect 12900 9392 12952 9444
rect 15108 9503 15160 9512
rect 15108 9469 15126 9503
rect 15126 9469 15160 9503
rect 15108 9460 15160 9469
rect 15384 9460 15436 9512
rect 18144 9528 18196 9580
rect 16396 9460 16448 9512
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 17684 9460 17736 9512
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 18512 9528 18564 9580
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 14924 9324 14976 9376
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 18788 9392 18840 9444
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 3148 9120 3200 9172
rect 4252 9120 4304 9172
rect 4712 9120 4764 9172
rect 2412 9052 2464 9104
rect 848 8959 900 8968
rect 848 8925 857 8959
rect 857 8925 891 8959
rect 891 8925 900 8959
rect 848 8916 900 8925
rect 1124 8959 1176 8968
rect 1124 8925 1133 8959
rect 1133 8925 1167 8959
rect 1167 8925 1176 8959
rect 1124 8916 1176 8925
rect 4160 8984 4212 9036
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 2596 8823 2648 8832
rect 2596 8789 2605 8823
rect 2605 8789 2639 8823
rect 2639 8789 2648 8823
rect 2596 8780 2648 8789
rect 2688 8780 2740 8832
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 4712 8916 4764 8968
rect 6184 9120 6236 9172
rect 6736 9052 6788 9104
rect 8852 9120 8904 9172
rect 9496 9120 9548 9172
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 9588 9052 9640 9104
rect 10416 9052 10468 9104
rect 10876 9052 10928 9104
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 8760 8984 8812 9036
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 8116 8916 8168 8968
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 3884 8780 3936 8832
rect 8300 8848 8352 8900
rect 4804 8780 4856 8832
rect 9772 8780 9824 8832
rect 10324 8984 10376 9036
rect 11520 9052 11572 9104
rect 11796 9163 11848 9172
rect 11796 9129 11805 9163
rect 11805 9129 11839 9163
rect 11839 9129 11848 9163
rect 11796 9120 11848 9129
rect 12808 9120 12860 9172
rect 14464 9120 14516 9172
rect 12164 9052 12216 9104
rect 13360 8984 13412 9036
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 15568 9095 15620 9104
rect 15568 9061 15577 9095
rect 15577 9061 15611 9095
rect 15611 9061 15620 9095
rect 15568 9052 15620 9061
rect 16396 9052 16448 9104
rect 10876 8916 10928 8968
rect 12716 8916 12768 8968
rect 14464 8916 14516 8968
rect 10784 8780 10836 8832
rect 11796 8848 11848 8900
rect 12164 8848 12216 8900
rect 15016 8984 15068 9036
rect 15108 8984 15160 9036
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 16764 8984 16816 9036
rect 17224 8984 17276 9036
rect 17868 8984 17920 9036
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 18420 8916 18472 8968
rect 16488 8848 16540 8900
rect 18604 8848 18656 8900
rect 13268 8780 13320 8832
rect 16120 8780 16172 8832
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 1124 8576 1176 8628
rect 3608 8576 3660 8628
rect 5356 8576 5408 8628
rect 4620 8508 4672 8560
rect 8760 8508 8812 8560
rect 9036 8576 9088 8628
rect 11152 8576 11204 8628
rect 11980 8576 12032 8628
rect 12072 8619 12124 8628
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 848 8440 900 8492
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 6828 8440 6880 8492
rect 8300 8440 8352 8492
rect 11060 8440 11112 8492
rect 1584 8372 1636 8424
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2596 8372 2648 8424
rect 5816 8372 5868 8424
rect 7288 8372 7340 8424
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 10324 8372 10376 8424
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 2504 8304 2556 8356
rect 1952 8236 2004 8288
rect 2412 8236 2464 8288
rect 6920 8304 6972 8356
rect 8024 8304 8076 8356
rect 10876 8304 10928 8356
rect 10968 8304 11020 8356
rect 11152 8304 11204 8356
rect 11888 8372 11940 8424
rect 12440 8372 12492 8424
rect 12164 8304 12216 8356
rect 12992 8372 13044 8424
rect 18328 8576 18380 8628
rect 16580 8508 16632 8560
rect 18420 8551 18472 8560
rect 14004 8440 14056 8492
rect 14740 8440 14792 8492
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 8760 8236 8812 8288
rect 11428 8236 11480 8288
rect 12440 8236 12492 8288
rect 12532 8279 12584 8288
rect 12532 8245 12541 8279
rect 12541 8245 12575 8279
rect 12575 8245 12584 8279
rect 12532 8236 12584 8245
rect 12992 8236 13044 8288
rect 14280 8372 14332 8424
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 17408 8440 17460 8492
rect 17776 8440 17828 8492
rect 18420 8517 18429 8551
rect 18429 8517 18463 8551
rect 18463 8517 18472 8551
rect 18420 8508 18472 8517
rect 18880 8508 18932 8560
rect 15108 8372 15160 8424
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 16212 8372 16264 8424
rect 16396 8372 16448 8424
rect 17592 8372 17644 8424
rect 15016 8304 15068 8356
rect 17868 8304 17920 8356
rect 15292 8236 15344 8288
rect 18236 8236 18288 8288
rect 18696 8279 18748 8288
rect 18696 8245 18705 8279
rect 18705 8245 18739 8279
rect 18739 8245 18748 8279
rect 18696 8236 18748 8245
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 1860 8075 1912 8084
rect 1860 8041 1869 8075
rect 1869 8041 1903 8075
rect 1903 8041 1912 8075
rect 1860 8032 1912 8041
rect 1952 8032 2004 8084
rect 7012 8032 7064 8084
rect 7380 8032 7432 8084
rect 7840 8032 7892 8084
rect 1584 7964 1636 8016
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 7196 7896 7248 7948
rect 8116 8007 8168 8016
rect 8116 7973 8125 8007
rect 8125 7973 8159 8007
rect 8159 7973 8168 8007
rect 8116 7964 8168 7973
rect 8484 8032 8536 8084
rect 8576 7964 8628 8016
rect 8760 8007 8812 8016
rect 8760 7973 8769 8007
rect 8769 7973 8803 8007
rect 8803 7973 8812 8007
rect 8760 7964 8812 7973
rect 10232 8032 10284 8084
rect 10784 7964 10836 8016
rect 11520 7964 11572 8016
rect 7288 7828 7340 7880
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 9404 7896 9456 7948
rect 9772 7896 9824 7948
rect 10508 7896 10560 7948
rect 11244 7896 11296 7948
rect 11704 7939 11756 7948
rect 11704 7905 11713 7939
rect 11713 7905 11747 7939
rect 11747 7905 11756 7939
rect 11704 7896 11756 7905
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 12440 7896 12492 7948
rect 12992 7896 13044 7948
rect 13176 7939 13228 7948
rect 13176 7905 13185 7939
rect 13185 7905 13219 7939
rect 13219 7905 13228 7939
rect 13176 7896 13228 7905
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 13728 7896 13780 7948
rect 15016 7896 15068 7948
rect 15108 7939 15160 7948
rect 15108 7905 15117 7939
rect 15117 7905 15151 7939
rect 15151 7905 15160 7939
rect 15108 7896 15160 7905
rect 10232 7828 10284 7880
rect 10416 7828 10468 7880
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 4068 7692 4120 7744
rect 12440 7760 12492 7812
rect 12624 7760 12676 7812
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 13636 7760 13688 7812
rect 14004 7760 14056 7812
rect 14372 7760 14424 7812
rect 14556 7803 14608 7812
rect 14556 7769 14565 7803
rect 14565 7769 14599 7803
rect 14599 7769 14608 7803
rect 14556 7760 14608 7769
rect 15016 7803 15068 7812
rect 15016 7769 15025 7803
rect 15025 7769 15059 7803
rect 15059 7769 15068 7803
rect 15016 7760 15068 7769
rect 18420 8032 18472 8084
rect 18604 8032 18656 8084
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 17592 7896 17644 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 18512 7939 18564 7948
rect 18512 7905 18521 7939
rect 18521 7905 18555 7939
rect 18555 7905 18564 7939
rect 18512 7896 18564 7905
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 17776 7760 17828 7812
rect 9680 7692 9732 7744
rect 10416 7692 10468 7744
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 11980 7692 12032 7744
rect 13084 7735 13136 7744
rect 13084 7701 13093 7735
rect 13093 7701 13127 7735
rect 13127 7701 13136 7735
rect 13084 7692 13136 7701
rect 13452 7692 13504 7744
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 2504 7488 2556 7540
rect 848 7395 900 7404
rect 848 7361 857 7395
rect 857 7361 891 7395
rect 891 7361 900 7395
rect 848 7352 900 7361
rect 2412 7284 2464 7336
rect 1124 7259 1176 7268
rect 1124 7225 1133 7259
rect 1133 7225 1167 7259
rect 1167 7225 1176 7259
rect 1124 7216 1176 7225
rect 5448 7488 5500 7540
rect 5816 7488 5868 7540
rect 10324 7488 10376 7540
rect 11704 7488 11756 7540
rect 7012 7420 7064 7472
rect 4160 7352 4212 7404
rect 6828 7352 6880 7404
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 2964 7216 3016 7268
rect 7564 7216 7616 7268
rect 3792 7191 3844 7200
rect 3792 7157 3801 7191
rect 3801 7157 3835 7191
rect 3835 7157 3844 7191
rect 3792 7148 3844 7157
rect 4252 7148 4304 7200
rect 6920 7148 6972 7200
rect 7380 7148 7432 7200
rect 8024 7284 8076 7336
rect 8116 7284 8168 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8852 7352 8904 7404
rect 9680 7352 9732 7404
rect 9312 7216 9364 7268
rect 9772 7284 9824 7336
rect 12532 7420 12584 7472
rect 10232 7284 10284 7336
rect 11336 7284 11388 7336
rect 11428 7327 11480 7336
rect 11428 7293 11437 7327
rect 11437 7293 11471 7327
rect 11471 7293 11480 7327
rect 11428 7284 11480 7293
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 11796 7284 11848 7336
rect 13360 7420 13412 7472
rect 13728 7463 13780 7472
rect 13728 7429 13737 7463
rect 13737 7429 13771 7463
rect 13771 7429 13780 7463
rect 13728 7420 13780 7429
rect 14096 7488 14148 7540
rect 18696 7488 18748 7540
rect 18880 7488 18932 7540
rect 14556 7420 14608 7472
rect 10232 7148 10284 7200
rect 10416 7148 10468 7200
rect 11152 7216 11204 7268
rect 12072 7259 12124 7268
rect 12072 7225 12081 7259
rect 12081 7225 12115 7259
rect 12115 7225 12124 7259
rect 12072 7216 12124 7225
rect 11060 7148 11112 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 11704 7148 11756 7200
rect 14096 7284 14148 7336
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 13268 7216 13320 7268
rect 18052 7420 18104 7472
rect 18144 7420 18196 7472
rect 18328 7420 18380 7472
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 17776 7352 17828 7404
rect 15844 7284 15896 7336
rect 16028 7284 16080 7336
rect 17684 7284 17736 7336
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 18236 7216 18288 7268
rect 13084 7148 13136 7200
rect 18696 7148 18748 7200
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 1952 6944 2004 6996
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 4068 6944 4120 6996
rect 4160 6944 4212 6996
rect 7196 6944 7248 6996
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 1124 6740 1176 6792
rect 5264 6876 5316 6928
rect 4344 6808 4396 6860
rect 5356 6808 5408 6860
rect 10416 6944 10468 6996
rect 10508 6944 10560 6996
rect 10048 6919 10100 6928
rect 10048 6885 10057 6919
rect 10057 6885 10091 6919
rect 10091 6885 10100 6919
rect 11612 6987 11664 6996
rect 11612 6953 11621 6987
rect 11621 6953 11655 6987
rect 11655 6953 11664 6987
rect 11612 6944 11664 6953
rect 10048 6876 10100 6885
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 4804 6672 4856 6724
rect 4988 6672 5040 6724
rect 2504 6604 2556 6656
rect 3792 6604 3844 6656
rect 4896 6604 4948 6656
rect 5448 6604 5500 6656
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 8300 6740 8352 6792
rect 8760 6740 8812 6792
rect 9680 6740 9732 6792
rect 11336 6808 11388 6860
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 7380 6604 7432 6656
rect 9404 6647 9456 6656
rect 9404 6613 9413 6647
rect 9413 6613 9447 6647
rect 9447 6613 9456 6647
rect 9404 6604 9456 6613
rect 10876 6604 10928 6656
rect 11796 6876 11848 6928
rect 11612 6808 11664 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 12900 6808 12952 6860
rect 15568 6944 15620 6996
rect 13820 6876 13872 6928
rect 14372 6876 14424 6928
rect 15200 6876 15252 6928
rect 15292 6808 15344 6860
rect 11888 6672 11940 6724
rect 12808 6672 12860 6724
rect 11612 6604 11664 6656
rect 11704 6604 11756 6656
rect 12348 6604 12400 6656
rect 13452 6672 13504 6724
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 14004 6740 14056 6792
rect 15108 6740 15160 6792
rect 15844 6851 15896 6860
rect 15844 6817 15853 6851
rect 15853 6817 15887 6851
rect 15887 6817 15896 6851
rect 15844 6808 15896 6817
rect 16764 6876 16816 6928
rect 17592 6876 17644 6928
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 15476 6740 15528 6792
rect 18144 6808 18196 6860
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 15384 6672 15436 6724
rect 15752 6672 15804 6724
rect 16028 6672 16080 6724
rect 16396 6715 16448 6724
rect 16396 6681 16405 6715
rect 16405 6681 16439 6715
rect 16439 6681 16448 6715
rect 16396 6672 16448 6681
rect 16764 6672 16816 6724
rect 17776 6740 17828 6792
rect 13176 6604 13228 6613
rect 15936 6604 15988 6656
rect 16580 6604 16632 6656
rect 16856 6604 16908 6656
rect 17224 6604 17276 6656
rect 17960 6604 18012 6656
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 3976 6400 4028 6452
rect 4344 6400 4396 6452
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 6092 6443 6144 6452
rect 6092 6409 6101 6443
rect 6101 6409 6135 6443
rect 6135 6409 6144 6443
rect 6092 6400 6144 6409
rect 6276 6400 6328 6452
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5264 6264 5316 6316
rect 3976 6128 4028 6180
rect 4068 6171 4120 6180
rect 4068 6137 4077 6171
rect 4077 6137 4111 6171
rect 4111 6137 4120 6171
rect 4068 6128 4120 6137
rect 4160 6128 4212 6180
rect 5080 6196 5132 6248
rect 4436 6103 4488 6112
rect 4436 6069 4445 6103
rect 4445 6069 4479 6103
rect 4479 6069 4488 6103
rect 4436 6060 4488 6069
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 13820 6400 13872 6452
rect 14188 6443 14240 6452
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 15660 6400 15712 6452
rect 17500 6400 17552 6452
rect 18236 6443 18288 6452
rect 18236 6409 18245 6443
rect 18245 6409 18279 6443
rect 18279 6409 18288 6443
rect 18236 6400 18288 6409
rect 8300 6264 8352 6316
rect 8392 6264 8444 6316
rect 5356 6128 5408 6180
rect 8484 6196 8536 6248
rect 11336 6332 11388 6384
rect 12624 6375 12676 6384
rect 12624 6341 12633 6375
rect 12633 6341 12667 6375
rect 12667 6341 12676 6375
rect 12624 6332 12676 6341
rect 9128 6264 9180 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 9404 6264 9456 6316
rect 10140 6264 10192 6316
rect 13176 6264 13228 6316
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16028 6264 16080 6316
rect 16764 6264 16816 6316
rect 10048 6128 10100 6180
rect 5448 6060 5500 6112
rect 6460 6060 6512 6112
rect 8300 6060 8352 6112
rect 8576 6060 8628 6112
rect 9496 6060 9548 6112
rect 10508 6128 10560 6180
rect 10876 6060 10928 6112
rect 12900 6196 12952 6248
rect 12532 6128 12584 6180
rect 12808 6171 12860 6180
rect 12808 6137 12817 6171
rect 12817 6137 12851 6171
rect 12851 6137 12860 6171
rect 12808 6128 12860 6137
rect 12992 6060 13044 6112
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 14372 6196 14424 6248
rect 14464 6196 14516 6248
rect 15844 6239 15896 6248
rect 13820 6128 13872 6180
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 18604 6332 18656 6384
rect 17500 6264 17552 6316
rect 18328 6264 18380 6316
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 17776 6239 17828 6248
rect 15752 6128 15804 6180
rect 16948 6128 17000 6180
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 17960 6239 18012 6248
rect 17960 6205 17969 6239
rect 17969 6205 18003 6239
rect 18003 6205 18012 6239
rect 17960 6196 18012 6205
rect 17592 6171 17644 6180
rect 17592 6137 17601 6171
rect 17601 6137 17635 6171
rect 17635 6137 17644 6171
rect 17592 6128 17644 6137
rect 17224 6060 17276 6112
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 18788 6196 18840 6248
rect 18420 6060 18472 6112
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 2412 5856 2464 5908
rect 2504 5831 2556 5840
rect 2504 5797 2513 5831
rect 2513 5797 2547 5831
rect 2547 5797 2556 5831
rect 2504 5788 2556 5797
rect 848 5720 900 5772
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 4344 5856 4396 5908
rect 4436 5856 4488 5908
rect 4804 5856 4856 5908
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 8576 5856 8628 5908
rect 9220 5856 9272 5908
rect 10876 5856 10928 5908
rect 9588 5788 9640 5840
rect 5540 5720 5592 5772
rect 7288 5763 7340 5772
rect 7288 5729 7297 5763
rect 7297 5729 7331 5763
rect 7331 5729 7340 5763
rect 7288 5720 7340 5729
rect 7380 5720 7432 5772
rect 4804 5584 4856 5636
rect 4988 5584 5040 5636
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6920 5652 6972 5704
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 4436 5516 4488 5568
rect 8300 5652 8352 5704
rect 9312 5584 9364 5636
rect 11520 5856 11572 5908
rect 11428 5788 11480 5840
rect 15476 5856 15528 5908
rect 15568 5856 15620 5908
rect 17684 5856 17736 5908
rect 10416 5652 10468 5704
rect 10968 5652 11020 5704
rect 11980 5720 12032 5772
rect 11796 5652 11848 5704
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 12716 5720 12768 5772
rect 13360 5652 13412 5704
rect 13636 5720 13688 5772
rect 14096 5720 14148 5772
rect 15384 5720 15436 5772
rect 18604 5831 18656 5840
rect 18604 5797 18613 5831
rect 18613 5797 18647 5831
rect 18647 5797 18656 5831
rect 18604 5788 18656 5797
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 15936 5720 15988 5772
rect 16396 5720 16448 5772
rect 17224 5763 17276 5772
rect 17224 5729 17233 5763
rect 17233 5729 17267 5763
rect 17267 5729 17276 5763
rect 17224 5720 17276 5729
rect 7932 5516 7984 5568
rect 12716 5516 12768 5568
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 13728 5516 13780 5568
rect 15752 5584 15804 5636
rect 15200 5516 15252 5568
rect 15292 5516 15344 5568
rect 16304 5652 16356 5704
rect 18512 5720 18564 5772
rect 18880 5763 18932 5772
rect 18880 5729 18889 5763
rect 18889 5729 18923 5763
rect 18923 5729 18932 5763
rect 18880 5720 18932 5729
rect 18052 5652 18104 5704
rect 18972 5652 19024 5704
rect 16948 5584 17000 5636
rect 18512 5584 18564 5636
rect 16120 5516 16172 5568
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 4160 5312 4212 5364
rect 3792 5176 3844 5228
rect 7196 5312 7248 5364
rect 5448 5176 5500 5228
rect 4804 5108 4856 5160
rect 6736 5244 6788 5296
rect 8392 5312 8444 5364
rect 8852 5312 8904 5364
rect 8116 5244 8168 5296
rect 10416 5312 10468 5364
rect 10600 5244 10652 5296
rect 6920 5108 6972 5160
rect 9404 5176 9456 5228
rect 9680 5176 9732 5228
rect 10784 5176 10836 5228
rect 10692 5108 10744 5160
rect 8024 5040 8076 5092
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 9312 5040 9364 5092
rect 9496 5040 9548 5092
rect 11060 5108 11112 5160
rect 12532 5312 12584 5364
rect 13360 5312 13412 5364
rect 16120 5355 16172 5364
rect 16120 5321 16129 5355
rect 16129 5321 16163 5355
rect 16163 5321 16172 5355
rect 16120 5312 16172 5321
rect 18420 5312 18472 5364
rect 11612 5244 11664 5296
rect 13820 5244 13872 5296
rect 14096 5244 14148 5296
rect 15660 5244 15712 5296
rect 15752 5287 15804 5296
rect 15752 5253 15761 5287
rect 15761 5253 15795 5287
rect 15795 5253 15804 5287
rect 15752 5244 15804 5253
rect 15844 5244 15896 5296
rect 16212 5244 16264 5296
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 12716 5176 12768 5228
rect 11980 5108 12032 5160
rect 12256 5151 12308 5160
rect 12256 5117 12265 5151
rect 12265 5117 12299 5151
rect 12299 5117 12308 5151
rect 12256 5108 12308 5117
rect 12992 5108 13044 5160
rect 9404 4972 9456 5024
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 11520 4972 11572 5024
rect 11980 4972 12032 5024
rect 12992 4972 13044 5024
rect 13360 4972 13412 5024
rect 15292 5108 15344 5160
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 16304 5108 16356 5117
rect 14004 5040 14056 5092
rect 15660 5040 15712 5092
rect 16580 5151 16632 5160
rect 16580 5117 16589 5151
rect 16589 5117 16623 5151
rect 16623 5117 16632 5151
rect 16580 5108 16632 5117
rect 16488 5040 16540 5092
rect 17500 5108 17552 5160
rect 17592 5108 17644 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 18972 5151 19024 5160
rect 18972 5117 18981 5151
rect 18981 5117 19015 5151
rect 19015 5117 19024 5151
rect 18972 5108 19024 5117
rect 17408 5040 17460 5092
rect 18052 5040 18104 5092
rect 14280 4972 14332 5024
rect 17224 4972 17276 5024
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 3792 4768 3844 4820
rect 480 4632 532 4684
rect 4436 4700 4488 4752
rect 4804 4700 4856 4752
rect 6460 4768 6512 4820
rect 7196 4768 7248 4820
rect 8024 4768 8076 4820
rect 10416 4768 10468 4820
rect 11428 4768 11480 4820
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 11796 4768 11848 4820
rect 12256 4768 12308 4820
rect 16120 4768 16172 4820
rect 16212 4811 16264 4820
rect 16212 4777 16221 4811
rect 16221 4777 16255 4811
rect 16255 4777 16264 4811
rect 16212 4768 16264 4777
rect 17408 4811 17460 4820
rect 17408 4777 17417 4811
rect 17417 4777 17451 4811
rect 17451 4777 17460 4811
rect 17408 4768 17460 4777
rect 17868 4768 17920 4820
rect 10968 4700 11020 4752
rect 12164 4700 12216 4752
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 7932 4564 7984 4616
rect 10232 4632 10284 4684
rect 11612 4632 11664 4684
rect 15384 4632 15436 4684
rect 16672 4700 16724 4752
rect 15936 4632 15988 4684
rect 16304 4632 16356 4684
rect 8852 4607 8904 4616
rect 8852 4573 8861 4607
rect 8861 4573 8895 4607
rect 8895 4573 8904 4607
rect 8852 4564 8904 4573
rect 9220 4564 9272 4616
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 11060 4564 11112 4616
rect 12532 4564 12584 4616
rect 13728 4564 13780 4616
rect 16488 4564 16540 4616
rect 17132 4675 17184 4684
rect 17132 4641 17141 4675
rect 17141 4641 17175 4675
rect 17175 4641 17184 4675
rect 17132 4632 17184 4641
rect 17316 4632 17368 4684
rect 19156 4632 19208 4684
rect 18052 4564 18104 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 14832 4496 14884 4548
rect 1032 4471 1084 4480
rect 1032 4437 1041 4471
rect 1041 4437 1075 4471
rect 1075 4437 1084 4471
rect 1032 4428 1084 4437
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 10416 4428 10468 4480
rect 10508 4428 10560 4480
rect 11152 4428 11204 4480
rect 12164 4428 12216 4480
rect 14924 4428 14976 4480
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 8300 4224 8352 4276
rect 12808 4224 12860 4276
rect 17776 4224 17828 4276
rect 9220 4156 9272 4208
rect 848 4088 900 4140
rect 1032 4020 1084 4072
rect 7288 4088 7340 4140
rect 8208 4088 8260 4140
rect 3792 4020 3844 4072
rect 7932 4020 7984 4072
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 10692 4156 10744 4208
rect 11060 4088 11112 4140
rect 11520 4088 11572 4140
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 3608 3952 3660 4004
rect 6552 3995 6604 4004
rect 6552 3961 6561 3995
rect 6561 3961 6595 3995
rect 6595 3961 6604 3995
rect 6552 3952 6604 3961
rect 7196 3952 7248 4004
rect 10232 4020 10284 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 4896 3884 4948 3936
rect 8116 3884 8168 3936
rect 9220 3884 9272 3936
rect 10508 3884 10560 3936
rect 11520 3884 11572 3936
rect 12624 4156 12676 4208
rect 14832 4156 14884 4208
rect 13728 4063 13780 4072
rect 13728 4029 13737 4063
rect 13737 4029 13771 4063
rect 13771 4029 13780 4063
rect 13728 4020 13780 4029
rect 14004 4088 14056 4140
rect 16672 4156 16724 4208
rect 18052 4156 18104 4208
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 17224 4020 17276 4072
rect 18696 4020 18748 4072
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 16212 3952 16264 4004
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 2780 3680 2832 3732
rect 3608 3680 3660 3732
rect 6552 3680 6604 3732
rect 8116 3680 8168 3732
rect 9680 3680 9732 3732
rect 11152 3680 11204 3732
rect 8576 3612 8628 3664
rect 10508 3612 10560 3664
rect 11336 3612 11388 3664
rect 13728 3680 13780 3732
rect 14924 3612 14976 3664
rect 16304 3680 16356 3732
rect 17500 3723 17552 3732
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 8852 3476 8904 3528
rect 10416 3544 10468 3596
rect 12532 3476 12584 3528
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 17592 3587 17644 3596
rect 17592 3553 17601 3587
rect 17601 3553 17635 3587
rect 17635 3553 17644 3587
rect 17592 3544 17644 3553
rect 18144 3544 18196 3596
rect 18604 3544 18656 3596
rect 10784 3451 10836 3460
rect 10784 3417 10793 3451
rect 10793 3417 10827 3451
rect 10827 3417 10836 3451
rect 10784 3408 10836 3417
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 7380 3136 7432 3188
rect 16212 3136 16264 3188
rect 16764 3136 16816 3188
rect 7840 3068 7892 3120
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 7196 2864 7248 2916
rect 8208 2975 8260 2984
rect 8208 2941 8217 2975
rect 8217 2941 8251 2975
rect 8251 2941 8260 2975
rect 8208 2932 8260 2941
rect 10232 3000 10284 3052
rect 11428 3043 11480 3052
rect 11428 3009 11437 3043
rect 11437 3009 11471 3043
rect 11471 3009 11480 3043
rect 11428 3000 11480 3009
rect 14924 3068 14976 3120
rect 11980 3000 12032 3052
rect 11520 2932 11572 2984
rect 10692 2864 10744 2916
rect 7748 2796 7800 2848
rect 11704 2864 11756 2916
rect 14096 2932 14148 2984
rect 16212 3000 16264 3052
rect 17224 3000 17276 3052
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 17960 2975 18012 2984
rect 17960 2941 17969 2975
rect 17969 2941 18003 2975
rect 18003 2941 18012 2975
rect 17960 2932 18012 2941
rect 19708 2932 19760 2984
rect 14464 2864 14516 2916
rect 17500 2864 17552 2916
rect 13912 2796 13964 2848
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 16580 2592 16632 2644
rect 6736 2524 6788 2576
rect 6828 2524 6880 2576
rect 6092 2499 6144 2508
rect 6092 2465 6101 2499
rect 6101 2465 6135 2499
rect 6135 2465 6144 2499
rect 6092 2456 6144 2465
rect 7012 2456 7064 2508
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 10324 2456 10376 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 13176 2456 13228 2508
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 15844 2456 15896 2508
rect 10692 2388 10744 2440
rect 11612 2388 11664 2440
rect 11980 2388 12032 2440
rect 14464 2320 14516 2372
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 6920 2295 6972 2304
rect 6920 2261 6929 2295
rect 6929 2261 6963 2295
rect 6963 2261 6972 2295
rect 6920 2252 6972 2261
rect 11520 2252 11572 2304
rect 15752 2388 15804 2440
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19616 2456 19668 2508
rect 18236 2388 18288 2440
rect 17868 2320 17920 2372
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 6828 2048 6880 2100
rect 6920 2048 6972 2100
rect 9404 2048 9456 2100
rect 11796 2048 11848 2100
rect 15016 2048 15068 2100
rect 848 1887 900 1896
rect 848 1853 857 1887
rect 857 1853 891 1887
rect 891 1853 900 1887
rect 848 1844 900 1853
rect 5724 1887 5776 1896
rect 5724 1853 5733 1887
rect 5733 1853 5767 1887
rect 5767 1853 5776 1887
rect 5724 1844 5776 1853
rect 5816 1887 5868 1896
rect 5816 1853 5825 1887
rect 5825 1853 5859 1887
rect 5859 1853 5868 1887
rect 5816 1844 5868 1853
rect 14188 1980 14240 2032
rect 16212 2023 16264 2032
rect 16212 1989 16221 2023
rect 16221 1989 16255 2023
rect 16255 1989 16264 2023
rect 16212 1980 16264 1989
rect 17868 1980 17920 2032
rect 7288 1844 7340 1896
rect 7380 1887 7432 1896
rect 7380 1853 7389 1887
rect 7389 1853 7423 1887
rect 7423 1853 7432 1887
rect 7380 1844 7432 1853
rect 7472 1887 7524 1896
rect 7472 1853 7481 1887
rect 7481 1853 7515 1887
rect 7515 1853 7524 1887
rect 7472 1844 7524 1853
rect 7932 1887 7984 1896
rect 7932 1853 7941 1887
rect 7941 1853 7975 1887
rect 7975 1853 7984 1887
rect 7932 1844 7984 1853
rect 8024 1887 8076 1896
rect 8024 1853 8033 1887
rect 8033 1853 8067 1887
rect 8067 1853 8076 1887
rect 8024 1844 8076 1853
rect 8668 1844 8720 1896
rect 11612 1955 11664 1964
rect 11612 1921 11621 1955
rect 11621 1921 11655 1955
rect 11655 1921 11664 1955
rect 11612 1912 11664 1921
rect 9036 1844 9088 1896
rect 9680 1844 9732 1896
rect 10876 1844 10928 1896
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 14096 1912 14148 1964
rect 16764 1912 16816 1964
rect 9404 1776 9456 1828
rect 10324 1776 10376 1828
rect 11980 1844 12032 1896
rect 6092 1708 6144 1760
rect 11704 1708 11756 1760
rect 11980 1708 12032 1760
rect 14464 1844 14516 1896
rect 15016 1844 15068 1896
rect 15844 1887 15896 1896
rect 15844 1853 15853 1887
rect 15853 1853 15887 1887
rect 15887 1853 15896 1887
rect 15844 1844 15896 1853
rect 17960 1887 18012 1896
rect 17960 1853 17969 1887
rect 17969 1853 18003 1887
rect 18003 1853 18012 1887
rect 17960 1844 18012 1853
rect 18880 1887 18932 1896
rect 18880 1853 18889 1887
rect 18889 1853 18923 1887
rect 18923 1853 18932 1887
rect 18880 1844 18932 1853
rect 18512 1708 18564 1760
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 5816 1504 5868 1556
rect 6092 1368 6144 1420
rect 6920 1504 6972 1556
rect 7472 1504 7524 1556
rect 7932 1504 7984 1556
rect 10416 1504 10468 1556
rect 7104 1436 7156 1488
rect 6920 1411 6972 1420
rect 6920 1377 6929 1411
rect 6929 1377 6963 1411
rect 6963 1377 6972 1411
rect 6920 1368 6972 1377
rect 7196 1411 7248 1420
rect 7196 1377 7205 1411
rect 7205 1377 7239 1411
rect 7239 1377 7248 1411
rect 7196 1368 7248 1377
rect 7288 1411 7340 1420
rect 7288 1377 7297 1411
rect 7297 1377 7331 1411
rect 7331 1377 7340 1411
rect 7288 1368 7340 1377
rect 8668 1411 8720 1420
rect 8668 1377 8677 1411
rect 8677 1377 8711 1411
rect 8711 1377 8720 1411
rect 8668 1368 8720 1377
rect 9680 1368 9732 1420
rect 7104 1300 7156 1352
rect 7840 1300 7892 1352
rect 10692 1343 10744 1352
rect 10692 1309 10701 1343
rect 10701 1309 10735 1343
rect 10735 1309 10744 1343
rect 11520 1411 11572 1420
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 11980 1436 12032 1488
rect 15752 1479 15804 1488
rect 15752 1445 15761 1479
rect 15761 1445 15795 1479
rect 15795 1445 15804 1479
rect 15752 1436 15804 1445
rect 18512 1479 18564 1488
rect 18512 1445 18521 1479
rect 18521 1445 18555 1479
rect 18555 1445 18564 1479
rect 18512 1436 18564 1445
rect 13636 1411 13688 1420
rect 13636 1377 13645 1411
rect 13645 1377 13679 1411
rect 13679 1377 13688 1411
rect 13636 1368 13688 1377
rect 10692 1300 10744 1309
rect 10876 1300 10928 1352
rect 12624 1300 12676 1352
rect 13452 1300 13504 1352
rect 7288 1232 7340 1284
rect 9036 1275 9088 1284
rect 9036 1241 9045 1275
rect 9045 1241 9079 1275
rect 9079 1241 9088 1275
rect 9036 1232 9088 1241
rect 15476 1411 15528 1420
rect 15476 1377 15485 1411
rect 15485 1377 15519 1411
rect 15519 1377 15528 1411
rect 15476 1368 15528 1377
rect 17500 1411 17552 1420
rect 17500 1377 17509 1411
rect 17509 1377 17543 1411
rect 17543 1377 17552 1411
rect 17500 1368 17552 1377
rect 18236 1411 18288 1420
rect 18236 1377 18245 1411
rect 18245 1377 18279 1411
rect 18279 1377 18288 1411
rect 18236 1368 18288 1377
rect 19616 1368 19668 1420
rect 16120 1300 16172 1352
rect 17868 1343 17920 1352
rect 17868 1309 17877 1343
rect 17877 1309 17911 1343
rect 17911 1309 17920 1343
rect 17868 1300 17920 1309
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 6092 960 6144 1012
rect 6920 960 6972 1012
rect 7196 960 7248 1012
rect 19064 1003 19116 1012
rect 19064 969 19073 1003
rect 19073 969 19107 1003
rect 19107 969 19116 1003
rect 19064 960 19116 969
rect 3976 799 4028 808
rect 3976 765 3985 799
rect 3985 765 4019 799
rect 4019 765 4028 799
rect 3976 756 4028 765
rect 5724 756 5776 808
rect 7104 824 7156 876
rect 7380 824 7432 876
rect 6552 799 6604 808
rect 6552 765 6561 799
rect 6561 765 6595 799
rect 6595 765 6604 799
rect 6552 756 6604 765
rect 9036 824 9088 876
rect 10876 824 10928 876
rect 8668 688 8720 740
rect 9404 756 9456 808
rect 13636 935 13688 944
rect 13636 901 13645 935
rect 13645 901 13679 935
rect 13679 901 13688 935
rect 13636 892 13688 901
rect 17868 892 17920 944
rect 13452 824 13504 876
rect 14924 824 14976 876
rect 16120 867 16172 876
rect 16120 833 16129 867
rect 16129 833 16163 867
rect 16163 833 16172 867
rect 16120 824 16172 833
rect 11980 756 12032 808
rect 15016 756 15068 808
rect 17500 799 17552 808
rect 17500 765 17509 799
rect 17509 765 17543 799
rect 17543 765 17552 799
rect 17500 756 17552 765
rect 7288 620 7340 672
rect 15476 620 15528 672
rect 18052 620 18104 672
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 3882 19600 3938 20000
rect 7746 19600 7802 20000
rect 8390 19600 8446 20000
rect 9034 19600 9090 20000
rect 9678 19600 9734 20000
rect 10322 19600 10378 20000
rect 10966 19600 11022 20000
rect 15474 19600 15530 20000
rect 16118 19600 16174 20000
rect 18050 19600 18106 20000
rect 3896 18970 3924 19600
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 7760 18902 7788 19600
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 848 18760 900 18766
rect 848 18702 900 18708
rect 860 18465 888 18702
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 846 18456 902 18465
rect 2755 18459 3063 18468
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 846 18391 902 18400
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 4896 17808 4948 17814
rect 3606 17776 3662 17785
rect 4896 17750 4948 17756
rect 3606 17711 3662 17720
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 3436 15978 3464 16390
rect 3528 16114 3556 17614
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 848 14952 900 14958
rect 848 14894 900 14900
rect 860 14278 888 14894
rect 1124 14884 1176 14890
rect 1124 14826 1176 14832
rect 1136 14618 1164 14826
rect 1124 14612 1176 14618
rect 1124 14554 1176 14560
rect 1872 14482 1900 15302
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 3160 15026 3188 15506
rect 3528 15162 3556 16050
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2424 14498 2452 14554
rect 2700 14498 2728 14826
rect 2884 14550 2912 14962
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2332 14482 2452 14498
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2320 14476 2452 14482
rect 2372 14470 2452 14476
rect 2516 14470 2728 14498
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2320 14418 2372 14424
rect 848 14272 900 14278
rect 848 14214 900 14220
rect 2056 13802 2084 14418
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 14074 2176 14350
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 2056 13326 2084 13738
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 848 12776 900 12782
rect 848 12718 900 12724
rect 860 11218 888 12718
rect 1688 12434 1716 13262
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12850 1808 13126
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1596 12406 1716 12434
rect 1492 11824 1544 11830
rect 1492 11766 1544 11772
rect 848 11212 900 11218
rect 848 11154 900 11160
rect 1124 11144 1176 11150
rect 1124 11086 1176 11092
rect 1136 10810 1164 11086
rect 1124 10804 1176 10810
rect 1124 10746 1176 10752
rect 1504 10606 1532 11766
rect 1596 11694 1624 12406
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1596 9382 1624 11630
rect 1688 11558 1716 12242
rect 1872 12170 1900 13194
rect 2148 12238 2176 13330
rect 2516 12714 2544 14470
rect 2700 14414 2728 14470
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2608 14074 2636 14350
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 3160 13938 3188 14758
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3436 13870 3464 14894
rect 3528 14618 3556 15098
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 2424 11694 2452 12174
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 10606 1716 11494
rect 2424 11014 2452 11630
rect 2516 11286 2544 12650
rect 2608 12102 2636 12922
rect 3160 12918 3188 13330
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12374 2728 12650
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3068 12434 3096 12582
rect 3068 12406 3188 12434
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 3068 12170 3096 12406
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 3160 11676 3188 12406
rect 3252 12356 3280 12582
rect 3436 12434 3464 13806
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12782 3556 13126
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3436 12406 3556 12434
rect 3424 12368 3476 12374
rect 3252 12328 3424 12356
rect 3424 12310 3476 12316
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3240 11688 3292 11694
rect 3160 11648 3240 11676
rect 3240 11630 3292 11636
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10674 2452 10950
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 9654 1716 10542
rect 2608 10198 2636 11494
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 3160 10810 3188 11086
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 1124 8968 1176 8974
rect 1124 8910 1176 8916
rect 860 8498 888 8910
rect 1136 8634 1164 8910
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 860 7410 888 8434
rect 1596 8430 1624 9318
rect 1688 8430 1716 9590
rect 2516 9518 2544 10066
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 3160 9518 3188 10202
rect 3252 10130 3280 11630
rect 3344 10742 3372 11766
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3528 10674 3556 12406
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3436 9674 3464 10406
rect 3528 9994 3556 10610
rect 3620 10198 3648 17711
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3896 17338 3924 17614
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3712 15502 3740 16594
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3988 15638 4016 16186
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3896 15162 3924 15574
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3988 15026 4016 15574
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 15178 4108 15370
rect 4080 15150 4200 15178
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3988 12782 4016 14962
rect 4172 14958 4200 15150
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4080 14618 4108 14894
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4172 14550 4200 14894
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4264 14346 4292 14894
rect 4356 14482 4384 15846
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 15162 4660 15438
rect 4908 15178 4936 17750
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5460 17270 5488 17682
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5460 17134 5488 17206
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 4988 16176 5040 16182
rect 4988 16118 5040 16124
rect 4724 15162 4936 15178
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4724 15156 4948 15162
rect 4724 15150 4896 15156
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4264 13870 4292 14282
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4264 13462 4292 13806
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3712 12442 3740 12718
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 12442 3832 12582
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3792 12436 3844 12442
rect 3988 12434 4016 12718
rect 3988 12406 4108 12434
rect 3792 12378 3844 12384
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3436 9646 3556 9674
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1596 8022 1624 8366
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1872 8090 1900 8298
rect 1964 8294 1992 9454
rect 3160 9178 3188 9454
rect 3528 9382 3556 9646
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2424 8294 2452 9046
rect 3528 8974 3556 9318
rect 3516 8968 3568 8974
rect 2516 8894 2728 8922
rect 3516 8910 3568 8916
rect 2516 8362 2544 8894
rect 2700 8838 2728 8894
rect 3896 8838 3924 9930
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 2608 8430 2636 8774
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 3620 8634 3648 8774
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 1964 8090 1992 8230
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 848 7404 900 7410
rect 848 7346 900 7352
rect 860 5778 888 7346
rect 1124 7268 1176 7274
rect 1124 7210 1176 7216
rect 1136 6798 1164 7210
rect 1688 6866 1716 7686
rect 1964 7002 1992 8026
rect 2424 7342 2452 8230
rect 2516 7546 2544 8298
rect 4080 7750 4108 12406
rect 4172 12102 4200 12786
rect 4356 12714 4384 14418
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4356 12434 4384 12650
rect 4540 12458 4568 13194
rect 4724 12968 4752 15150
rect 4896 15098 4948 15104
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4816 14074 4844 15030
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4908 14618 4936 14894
rect 5000 14890 5028 16118
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 5460 15706 5488 17070
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5552 16658 5580 17002
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5644 16538 5672 17002
rect 5736 16998 5764 17682
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5828 17338 5856 17478
rect 6104 17338 6132 18090
rect 6380 17678 6408 18158
rect 8128 18086 8156 18770
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6840 17542 6868 18022
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6380 17270 6408 17478
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 6276 17128 6328 17134
rect 6380 17116 6408 17206
rect 6328 17088 6408 17116
rect 6644 17128 6696 17134
rect 6276 17070 6328 17076
rect 6644 17070 6696 17076
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 6656 16794 6684 17070
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 5552 16510 5672 16538
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5552 16454 5580 16510
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 14890 5212 15302
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 5000 14482 5028 14826
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 5460 14618 5488 15642
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4816 12986 4844 14010
rect 5000 13530 5028 14418
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4632 12940 4752 12968
rect 4804 12980 4856 12986
rect 4632 12764 4660 12940
rect 4804 12922 4856 12928
rect 4632 12736 4844 12764
rect 4356 12406 4476 12434
rect 4540 12430 4752 12458
rect 4448 12306 4476 12406
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11354 4200 12038
rect 4448 11558 4476 12242
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4172 10674 4200 11290
rect 4448 11286 4476 11494
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4632 11082 4660 11562
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4264 9178 4292 9318
rect 4724 9178 4752 12430
rect 4816 11898 4844 12736
rect 4908 12442 4936 13262
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 5000 12850 5028 13126
rect 5184 12986 5212 13330
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5276 12646 5304 12786
rect 5368 12646 5396 13398
rect 5460 13190 5488 14418
rect 5552 13938 5580 16390
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5736 15638 5764 15846
rect 5920 15706 5948 16526
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 5644 14550 5672 15506
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5920 14278 5948 15438
rect 6012 14550 6040 15506
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 6012 14074 6040 14486
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 6012 13530 6040 14010
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6104 13394 6132 15506
rect 6196 14346 6224 16594
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 15638 6408 16390
rect 6656 16250 6684 16730
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6748 15502 6776 16594
rect 6840 16454 6868 17478
rect 7116 17202 7144 17750
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7208 16998 7236 17478
rect 7300 17134 7328 17818
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7392 17338 7420 17750
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7116 16794 7144 16934
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 4896 12436 4948 12442
rect 6196 12434 6224 14282
rect 6564 13802 6592 15302
rect 6748 15162 6776 15438
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 14550 6776 14962
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 4896 12378 4948 12384
rect 6104 12406 6224 12434
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 10538 4844 11494
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1124 6792 1176 6798
rect 1124 6734 1176 6740
rect 2424 5914 2452 7278
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2976 6866 3004 7210
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3804 6662 3832 7142
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2516 5846 2544 6598
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 3988 6458 4016 7278
rect 4080 7002 4108 7686
rect 4172 7410 4200 8978
rect 4632 8566 4660 8978
rect 4712 8968 4764 8974
rect 4764 8928 4844 8956
rect 4712 8910 4764 8916
rect 4816 8838 4844 8928
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 7002 4200 7346
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3988 6186 4016 6394
rect 4172 6186 4200 6938
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 3988 5914 4016 6122
rect 4080 6066 4108 6122
rect 4264 6066 4292 7142
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6458 4384 6802
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4342 6352 4398 6361
rect 4342 6287 4398 6296
rect 4080 6038 4292 6066
rect 4356 5914 4384 6287
rect 4618 6216 4674 6225
rect 4618 6151 4674 6160
rect 4632 6118 4660 6151
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4448 5914 4476 6054
rect 4816 5914 4844 6666
rect 4908 6662 4936 11630
rect 5000 11354 5028 11630
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 5460 11354 5488 11494
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5460 11014 5488 11290
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5828 10674 5856 11698
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10810 6040 11154
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 5828 9586 5856 10610
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8634 5396 8978
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5828 8430 5856 8910
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 5828 7954 5856 8366
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5460 7546 5488 7890
rect 5828 7546 5856 7890
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 848 5772 900 5778
rect 848 5714 900 5720
rect 480 4684 532 4690
rect 480 4626 532 4632
rect 492 4185 520 4626
rect 478 4176 534 4185
rect 860 4146 888 5714
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 4172 5370 4200 5510
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4826 3832 5170
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 1032 4480 1084 4486
rect 1032 4422 1084 4428
rect 478 4111 534 4120
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 1044 4078 1072 4422
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 3804 4078 3832 4762
rect 4448 4758 4476 5510
rect 4816 5166 4844 5578
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4816 4758 4844 5102
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 1032 4072 1084 4078
rect 1032 4014 1084 4020
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3738 2820 3878
rect 3620 3738 3648 3946
rect 4908 3942 4936 6598
rect 5000 6458 5028 6666
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5170 6352 5226 6361
rect 5276 6322 5304 6870
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5170 6287 5172 6296
rect 5224 6287 5226 6296
rect 5264 6316 5316 6322
rect 5172 6258 5224 6264
rect 5264 6258 5316 6264
rect 5080 6248 5132 6254
rect 5000 6208 5080 6236
rect 5000 5642 5028 6208
rect 5080 6190 5132 6196
rect 5368 6186 5396 6802
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6338 5488 6598
rect 6104 6458 6132 12406
rect 6656 12306 6684 13874
rect 6748 13462 6776 14486
rect 6840 13734 6868 16390
rect 6932 16250 6960 16662
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6840 13326 6868 13670
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11762 6224 12038
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6472 11354 6500 12242
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6564 11286 6592 11562
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6564 10606 6592 11222
rect 6840 11150 6868 12786
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9586 6408 9862
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6196 8498 6224 9114
rect 6748 9110 6776 9386
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6458 6316 6734
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5460 6310 5580 6338
rect 5446 6216 5502 6225
rect 5356 6180 5408 6186
rect 5446 6151 5502 6160
rect 5356 6122 5408 6128
rect 5460 6118 5488 6151
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5460 5234 5488 6054
rect 5552 5778 5580 6310
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 6472 5710 6500 6054
rect 6748 5914 6776 9046
rect 6840 8498 6868 11086
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6840 7410 6868 8434
rect 6932 8362 6960 14894
rect 7024 14618 7052 15098
rect 7116 14822 7144 16730
rect 7208 16726 7236 16934
rect 7392 16726 7420 16934
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7208 14634 7236 16662
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 14606 7236 14634
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7024 13870 7052 14418
rect 7116 13870 7144 14606
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7024 9926 7052 13806
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13462 7144 13670
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7208 12986 7236 13806
rect 7300 13462 7328 14826
rect 7392 14006 7420 16662
rect 7576 16454 7604 17002
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7852 15366 7880 15846
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 7944 14618 7972 15506
rect 8220 15162 8248 15574
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8312 14958 8340 15846
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7484 13530 7512 13806
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7852 12850 7880 13942
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12918 8156 13126
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 11218 7236 12718
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12306 7880 12582
rect 8220 12442 8248 13262
rect 8312 13161 8340 13330
rect 8298 13152 8354 13161
rect 8298 13087 8354 13096
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8022 12336 8078 12345
rect 7472 12300 7524 12306
rect 7392 12260 7472 12288
rect 7392 11286 7420 12260
rect 7472 12242 7524 12248
rect 7840 12300 7892 12306
rect 8022 12271 8024 12280
rect 7840 12242 7892 12248
rect 8076 12271 8078 12280
rect 8116 12300 8168 12306
rect 8024 12242 8076 12248
rect 8116 12242 8168 12248
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7576 11354 7604 11834
rect 8128 11558 8156 12242
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 8312 11218 8340 13087
rect 8404 11286 8432 19600
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8496 15094 8524 15846
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 8496 12782 8524 15030
rect 8680 13394 8708 18634
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8956 17746 8984 18090
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8864 17134 8892 17614
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8772 16794 8800 17070
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8864 16114 8892 17070
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8864 14940 8892 16050
rect 8956 15638 8984 17682
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 8956 15502 8984 15574
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 15094 8984 15438
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8944 14952 8996 14958
rect 8864 14912 8944 14940
rect 8944 14894 8996 14900
rect 8956 14618 8984 14894
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8942 13424 8998 13433
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8864 13382 8942 13410
rect 8680 12986 8708 13330
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12434 8616 12718
rect 8496 12406 8616 12434
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7300 9382 7328 10134
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8430 7328 9318
rect 7838 8936 7894 8945
rect 7838 8871 7894 8880
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 7852 8430 7880 8871
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6932 7206 6960 8298
rect 7852 8090 7880 8366
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7024 7478 7052 8026
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7208 7002 7236 7890
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6748 5302 6776 5850
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 6932 5166 6960 5646
rect 7208 5370 7236 6938
rect 7300 5778 7328 7822
rect 7392 7206 7420 8026
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 7564 7268 7616 7274
rect 7944 7256 7972 9862
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8036 7342 8064 8298
rect 8128 8022 8156 8910
rect 8312 8906 8340 11154
rect 8390 10704 8446 10713
rect 8390 10639 8392 10648
rect 8444 10639 8446 10648
rect 8392 10610 8444 10616
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8404 9722 8432 10066
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8312 8498 8340 8842
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7426 8156 7958
rect 8128 7398 8248 7426
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 7616 7228 7972 7256
rect 7564 7210 7616 7216
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7944 6866 7972 7228
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 5778 7420 6598
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 6472 4826 6500 4966
rect 7208 4826 7236 5306
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7208 4010 7236 4762
rect 7288 4140 7340 4146
rect 7392 4128 7420 5714
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 7944 4622 7972 5510
rect 8036 5098 8064 7278
rect 8128 5302 8156 7278
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4826 8064 5034
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 7340 4100 7420 4128
rect 7288 4082 7340 4088
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 6564 3738 6592 3946
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 7392 3194 7420 4100
rect 7944 4078 7972 4558
rect 8220 4146 8248 7398
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 6322 8340 6734
rect 8404 6322 8432 9454
rect 8496 8090 8524 12406
rect 8680 11694 8708 12922
rect 8864 12850 8892 13382
rect 8942 13359 8998 13368
rect 8942 13288 8998 13297
rect 8942 13223 8944 13232
rect 8996 13223 8998 13232
rect 8944 13194 8996 13200
rect 8956 12850 8984 13194
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8758 12744 8814 12753
rect 9048 12730 9076 19600
rect 9692 18766 9720 19600
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9140 16590 9168 18702
rect 9220 18080 9272 18086
rect 9324 18068 9352 18702
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9272 18040 9352 18068
rect 9220 18022 9272 18028
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16114 9168 16526
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15706 9168 16050
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9232 15502 9260 15846
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13462 9168 13738
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 8758 12679 8814 12688
rect 8956 12702 9076 12730
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11354 8708 11630
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10606 8616 11018
rect 8680 10606 8708 11290
rect 8772 10742 8800 12679
rect 8956 12356 8984 12702
rect 9140 12646 9168 13398
rect 9232 12782 9260 15438
rect 9324 13512 9352 18040
rect 9692 17882 9720 18566
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 9827 17980 10135 17989
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 10244 17882 10272 18090
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16794 9720 16934
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15706 9628 15982
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 9600 15337 9628 15506
rect 9586 15328 9642 15337
rect 9586 15263 9642 15272
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9416 14618 9444 14826
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9692 14074 9720 14418
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9784 13870 9812 14010
rect 10152 13938 10180 14282
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10244 13870 10272 15506
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 9324 13484 9720 13512
rect 9324 13190 9352 13484
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9508 12918 9536 13330
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9416 12782 9444 12854
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9036 12368 9088 12374
rect 8956 12328 9036 12356
rect 9128 12368 9180 12374
rect 9036 12310 9088 12316
rect 9126 12336 9128 12345
rect 9180 12336 9182 12345
rect 9232 12306 9260 12718
rect 9126 12271 9182 12280
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9324 12170 9352 12718
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9312 12164 9364 12170
rect 9364 12124 9444 12152
rect 9312 12106 9364 12112
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11354 8892 11494
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 9586 8800 10406
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 9042 8800 9318
rect 8864 9178 8892 10542
rect 8956 10470 8984 11562
rect 9140 11558 9168 12106
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8772 8566 8800 8978
rect 9048 8634 9076 11290
rect 9140 11150 9168 11494
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9126 10976 9182 10985
rect 9126 10911 9182 10920
rect 9140 9586 9168 10911
rect 9232 10130 9260 12038
rect 9416 11762 9444 12124
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9324 10810 9352 11630
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11354 9444 11494
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9324 9586 9352 10746
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 9140 8430 9168 9318
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8772 8022 8800 8230
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5710 8340 6054
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8404 5370 8432 6258
rect 8496 6254 8524 7890
rect 8588 7342 8616 7958
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8772 6798 8800 7958
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7410 8892 7890
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 9140 6322 9168 8366
rect 9416 7954 9444 10746
rect 9508 10112 9536 12582
rect 9600 11082 9628 12582
rect 9692 12434 9720 13484
rect 10048 13320 10100 13326
rect 9862 13288 9918 13297
rect 10048 13262 10100 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9862 13223 9864 13232
rect 9916 13223 9918 13232
rect 9864 13194 9916 13200
rect 10060 12850 10088 13262
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9784 12646 9812 12786
rect 10244 12753 10272 13262
rect 10336 12986 10364 19600
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10230 12744 10286 12753
rect 10230 12679 10286 12688
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 9692 12406 9812 12434
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11354 9720 12106
rect 9784 11762 9812 12406
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11762 10088 12242
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11665 10088 11698
rect 10046 11656 10102 11665
rect 10046 11591 10102 11600
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 10244 11354 10272 12679
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10046 11248 10102 11257
rect 10046 11183 10048 11192
rect 10100 11183 10102 11192
rect 10232 11212 10284 11218
rect 10048 11154 10100 11160
rect 10336 11200 10364 12038
rect 10428 11898 10456 18702
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10520 17678 10548 18226
rect 10980 17898 11008 19600
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 15488 18834 15516 19600
rect 16132 18834 16160 19600
rect 18064 18834 18092 19600
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 10796 17870 11008 17898
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10520 17202 10548 17614
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10612 14396 10640 16934
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10704 14822 10732 15914
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10520 14368 10640 14396
rect 10520 13326 10548 14368
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13870 10640 14214
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10284 11172 10364 11200
rect 10232 11154 10284 11160
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9876 10674 9904 10950
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9968 10470 9996 11086
rect 10244 11082 10272 11154
rect 10232 11076 10284 11082
rect 10428 11064 10456 11222
rect 10232 11018 10284 11024
rect 10336 11036 10456 11064
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10742 10180 10950
rect 10140 10736 10192 10742
rect 10046 10704 10102 10713
rect 10140 10678 10192 10684
rect 10046 10639 10048 10648
rect 10100 10639 10102 10648
rect 10048 10610 10100 10616
rect 10152 10554 10180 10678
rect 10152 10526 10272 10554
rect 10336 10538 10364 11036
rect 10520 10996 10548 12582
rect 10612 12442 10640 13806
rect 10704 13462 10732 14282
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10704 12918 10732 13398
rect 10796 13326 10824 17870
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10980 17338 11008 17682
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 16114 11744 17138
rect 11900 16998 11928 17478
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 12544 17066 12572 17750
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17134 12664 17478
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14346 10916 14758
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13394 10916 13670
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10784 13320 10836 13326
rect 10980 13274 11008 14010
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10784 13262 10836 13268
rect 10888 13246 11008 13274
rect 10888 12918 10916 13246
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10692 12912 10744 12918
rect 10876 12912 10928 12918
rect 10692 12854 10744 12860
rect 10782 12880 10838 12889
rect 10876 12854 10928 12860
rect 10782 12815 10784 12824
rect 10836 12815 10838 12824
rect 10784 12786 10836 12792
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10690 12200 10746 12209
rect 10690 12135 10746 12144
rect 10704 11286 10732 12135
rect 10796 12102 10824 12650
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11286 10824 11494
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10428 10968 10548 10996
rect 9956 10464 10008 10470
rect 9692 10424 9956 10452
rect 9588 10124 9640 10130
rect 9508 10084 9588 10112
rect 9588 10066 9640 10072
rect 9692 10044 9720 10424
rect 9956 10406 10008 10412
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9692 10016 9904 10044
rect 9770 9888 9826 9897
rect 9770 9823 9826 9832
rect 9784 9704 9812 9823
rect 9876 9722 9904 10016
rect 9692 9676 9812 9704
rect 9864 9716 9916 9722
rect 9692 9568 9720 9676
rect 9864 9658 9916 9664
rect 9968 9674 9996 10202
rect 10244 10130 10272 10526
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10138 10024 10194 10033
rect 10060 9897 10088 9998
rect 10138 9959 10140 9968
rect 10192 9959 10194 9968
rect 10232 9988 10284 9994
rect 10140 9930 10192 9936
rect 10232 9930 10284 9936
rect 10046 9888 10102 9897
rect 10046 9823 10102 9832
rect 10244 9761 10272 9930
rect 10230 9752 10286 9761
rect 10230 9687 10286 9696
rect 9968 9646 10180 9674
rect 9600 9540 9720 9568
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 9178 9536 9454
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9600 9110 9628 9540
rect 10152 9518 10180 9646
rect 10140 9512 10192 9518
rect 10138 9480 10140 9489
rect 10232 9512 10284 9518
rect 10192 9480 10194 9489
rect 9680 9444 9732 9450
rect 10232 9454 10284 9460
rect 10138 9415 10194 9424
rect 9680 9386 9732 9392
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9692 7750 9720 9386
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 9862 8936 9918 8945
rect 9862 8871 9918 8880
rect 9772 8832 9824 8838
rect 9876 8820 9904 8871
rect 9824 8792 9904 8820
rect 9772 8774 9824 8780
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 10244 8090 10272 9454
rect 10336 9042 10364 10066
rect 10428 9518 10456 10968
rect 10612 10690 10640 11018
rect 10520 10662 10640 10690
rect 10520 9518 10548 10662
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 9722 10640 10134
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10704 9654 10732 11018
rect 10796 11014 10824 11222
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9324 6322 9352 7210
rect 9692 6798 9720 7346
rect 9784 7342 9812 7890
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10244 7342 10272 7822
rect 10336 7546 10364 8366
rect 10428 7886 10456 9046
rect 10506 8936 10562 8945
rect 10506 8871 10562 8880
rect 10520 7954 10548 8871
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10416 7880 10468 7886
rect 10468 7828 10548 7834
rect 10416 7822 10548 7828
rect 10428 7806 10548 7822
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10428 7206 10456 7686
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 6322 9444 6598
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 9140 5930 9168 6258
rect 9140 5914 9260 5930
rect 8576 5908 8628 5914
rect 9140 5908 9272 5914
rect 9140 5902 9220 5908
rect 8576 5850 8628 5856
rect 9220 5850 9272 5856
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4282 8340 4626
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8496 4185 8524 4422
rect 8482 4176 8538 4185
rect 8208 4140 8260 4146
rect 8482 4111 8538 4120
rect 8208 4082 8260 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3738 8156 3878
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8588 3670 8616 5850
rect 9324 5760 9352 6258
rect 9232 5732 9352 5760
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8864 4622 8892 5306
rect 9232 4622 9260 5732
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9324 5098 9352 5578
rect 9416 5234 9444 6258
rect 10060 6186 10088 6870
rect 10244 6338 10272 7142
rect 10428 7002 10456 7142
rect 10520 7002 10548 7806
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10152 6322 10272 6338
rect 10140 6316 10272 6322
rect 10192 6310 10272 6316
rect 10140 6258 10192 6264
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9508 5098 9536 6054
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9404 5024 9456 5030
rect 9600 4978 9628 5782
rect 10428 5710 10456 6938
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10428 5370 10456 5646
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9456 4972 9628 4978
rect 9404 4966 9628 4972
rect 9416 4950 9628 4966
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8864 3534 8892 4558
rect 9232 4214 9260 4558
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 9232 3942 9260 4150
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6840 2774 6868 2926
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 6748 2746 6868 2774
rect 6748 2582 6776 2746
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 848 1896 900 1902
rect 848 1838 900 1844
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 860 1465 888 1838
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 846 1456 902 1465
rect 846 1391 902 1400
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 5736 814 5764 1838
rect 5828 1562 5856 1838
rect 6104 1766 6132 2450
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6092 1760 6144 1766
rect 6092 1702 6144 1708
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 6104 1426 6132 1702
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6104 1018 6132 1158
rect 6092 1012 6144 1018
rect 6092 954 6144 960
rect 6564 814 6592 2246
rect 6840 2106 6868 2518
rect 7024 2514 7052 2926
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6920 2304 6972 2310
rect 7208 2258 7236 2858
rect 6920 2246 6972 2252
rect 6932 2106 6960 2246
rect 7024 2230 7236 2258
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 7024 1986 7052 2230
rect 7300 2122 7328 2926
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2514 7788 2790
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 6932 1958 7052 1986
rect 7116 2094 7328 2122
rect 6932 1562 6960 1958
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 7116 1494 7144 2094
rect 7288 1896 7340 1902
rect 7288 1838 7340 1844
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7472 1896 7524 1902
rect 7472 1838 7524 1844
rect 7104 1488 7156 1494
rect 7104 1430 7156 1436
rect 7300 1426 7328 1838
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 7196 1420 7248 1426
rect 7196 1362 7248 1368
rect 7288 1420 7340 1426
rect 7288 1362 7340 1368
rect 6932 1018 6960 1362
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 6920 1012 6972 1018
rect 6920 954 6972 960
rect 7116 882 7144 1294
rect 7208 1018 7236 1362
rect 7300 1290 7328 1362
rect 7288 1284 7340 1290
rect 7288 1226 7340 1232
rect 7196 1012 7248 1018
rect 7196 954 7248 960
rect 7104 876 7156 882
rect 7104 818 7156 824
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 5724 808 5776 814
rect 5724 750 5776 756
rect 6552 808 6604 814
rect 6552 750 6604 756
rect 3988 490 4016 750
rect 7300 678 7328 1226
rect 7392 882 7420 1838
rect 7484 1562 7512 1838
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7852 1358 7880 3062
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8220 2394 8248 2926
rect 8036 2366 8248 2394
rect 8036 1902 8064 2366
rect 9416 2106 9444 4558
rect 9600 4078 9628 4950
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9692 3738 9720 5170
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 10428 4826 10456 5306
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10244 4162 10272 4626
rect 10520 4486 10548 6122
rect 10612 5302 10640 9522
rect 10796 8838 10824 10542
rect 10888 10538 10916 12854
rect 10980 11234 11008 13126
rect 11072 12782 11100 13942
rect 11256 13870 11284 15642
rect 11440 15570 11468 16050
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11440 14958 11468 15506
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 11348 14618 11376 14894
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11256 13394 11284 13806
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11060 12368 11112 12374
rect 11058 12336 11060 12345
rect 11112 12336 11114 12345
rect 11058 12271 11114 12280
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11694 11100 12106
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11072 11354 11100 11630
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10980 11206 11100 11234
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10888 10130 10916 10474
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9518 10916 10066
rect 11072 9926 11100 11206
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10980 9722 11008 9862
rect 11058 9752 11114 9761
rect 10968 9716 11020 9722
rect 11058 9687 11114 9696
rect 10968 9658 11020 9664
rect 11072 9518 11100 9687
rect 11164 9586 11192 13330
rect 11348 12986 11376 13670
rect 11440 13161 11468 13738
rect 11532 13394 11560 15914
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15706 11652 15846
rect 11716 15706 11744 16050
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11716 14414 11744 15642
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11900 13394 11928 16934
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15706 12112 15982
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11426 13152 11482 13161
rect 11426 13087 11482 13096
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11256 11694 11284 12310
rect 11440 12306 11468 13087
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11532 11778 11560 12718
rect 11624 12442 11652 12922
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11610 12336 11666 12345
rect 11716 12322 11744 13330
rect 11992 13274 12020 14418
rect 11666 12294 11744 12322
rect 11900 13246 12020 13274
rect 11796 12300 11848 12306
rect 11610 12271 11666 12280
rect 11796 12242 11848 12248
rect 11348 11750 11560 11778
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11348 10742 11376 11750
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11704 11688 11756 11694
rect 11808 11676 11836 12242
rect 11756 11648 11836 11676
rect 11704 11630 11756 11636
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 10130 11284 10406
rect 11348 10266 11376 10678
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11348 9674 11376 10202
rect 11440 9761 11468 11630
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11218 11560 11562
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11716 11150 11744 11630
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11624 10810 11652 11018
rect 11716 10962 11744 11086
rect 11716 10934 11836 10962
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11426 9752 11482 9761
rect 11426 9687 11482 9696
rect 11256 9646 11376 9674
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10876 9512 10928 9518
rect 11060 9512 11112 9518
rect 10876 9454 10928 9460
rect 10966 9480 11022 9489
rect 11060 9454 11112 9460
rect 11150 9480 11206 9489
rect 10966 9415 11022 9424
rect 11150 9415 11206 9424
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10888 8974 10916 9046
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8022 10824 8774
rect 10888 8362 10916 8910
rect 10980 8362 11008 9415
rect 11164 8634 11192 9415
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11150 8528 11206 8537
rect 11060 8492 11112 8498
rect 11150 8463 11206 8472
rect 11060 8434 11112 8440
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 11072 7206 11100 8434
rect 11164 8362 11192 8463
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11256 7954 11284 9646
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11348 9178 11376 9454
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11440 8378 11468 9522
rect 11532 9110 11560 10066
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11348 8350 11468 8378
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11164 6798 11192 7210
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6118 10916 6598
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5914 10916 6054
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10244 4134 10364 4162
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 10244 3058 10272 4014
rect 10336 3482 10364 4134
rect 10428 3602 10456 4422
rect 10704 4214 10732 5102
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3670 10548 3878
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10336 3454 10456 3482
rect 10796 3466 10824 5170
rect 10980 4758 11008 5646
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11072 4622 11100 5102
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4146 11100 4558
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11164 3738 11192 4422
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10232 3052 10284 3058
rect 10284 3012 10364 3040
rect 10232 2994 10284 3000
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 10336 2514 10364 3012
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 7932 1896 7984 1902
rect 7932 1838 7984 1844
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 7944 1562 7972 1838
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8680 1426 8708 1838
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 7380 876 7432 882
rect 7380 818 7432 824
rect 8680 746 8708 1362
rect 9048 1290 9076 1838
rect 9404 1828 9456 1834
rect 9404 1770 9456 1776
rect 9036 1284 9088 1290
rect 9036 1226 9088 1232
rect 9048 882 9076 1226
rect 9036 876 9088 882
rect 9036 818 9088 824
rect 9416 814 9444 1770
rect 9692 1426 9720 1838
rect 10336 1834 10364 2450
rect 10324 1828 10376 1834
rect 10324 1770 10376 1776
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 10428 1562 10456 3454
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10704 2446 10732 2858
rect 11256 2774 11284 7686
rect 11348 7342 11376 8350
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 7342 11468 8230
rect 11532 8129 11560 8366
rect 11518 8120 11574 8129
rect 11518 8055 11574 8064
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11348 6866 11376 7278
rect 11532 7206 11560 7958
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11348 6390 11376 6802
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11426 5944 11482 5953
rect 11532 5914 11560 7142
rect 11624 7002 11652 9386
rect 11716 8265 11744 9862
rect 11808 9466 11836 10934
rect 11900 9586 11928 13246
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11808 9438 11928 9466
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11808 9178 11836 9318
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11702 8256 11758 8265
rect 11702 8191 11758 8200
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7546 11744 7890
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11702 7440 11758 7449
rect 11702 7375 11758 7384
rect 11716 7342 11744 7375
rect 11808 7342 11836 8842
rect 11900 8514 11928 9438
rect 11992 8634 12020 13126
rect 12084 12968 12112 15642
rect 12268 15638 12296 15846
rect 12544 15638 12572 17002
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 12532 15632 12584 15638
rect 12532 15574 12584 15580
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 12544 15026 12572 15574
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12360 13530 12388 13738
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12162 13424 12218 13433
rect 12544 13394 12572 14350
rect 12636 13870 12664 17070
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 14482 13400 14758
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12162 13359 12164 13368
rect 12216 13359 12218 13368
rect 12532 13388 12584 13394
rect 12164 13330 12216 13336
rect 12532 13330 12584 13336
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 12544 12986 12572 13126
rect 12728 12986 12756 13126
rect 12532 12980 12584 12986
rect 12084 12940 12204 12968
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 8634 12112 12582
rect 12176 12374 12204 12940
rect 12532 12922 12584 12928
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12254 12336 12310 12345
rect 12360 12306 12388 12854
rect 12820 12782 12848 13670
rect 12912 13394 12940 14282
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13394 13032 14214
rect 13096 13394 13124 14418
rect 14936 13870 14964 14554
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 15028 14006 15056 14486
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13372 13394 13400 13738
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12254 12271 12310 12280
rect 12348 12300 12400 12306
rect 12268 12170 12296 12271
rect 12348 12242 12400 12248
rect 12360 12209 12388 12242
rect 12346 12200 12402 12209
rect 12256 12164 12308 12170
rect 12346 12135 12402 12144
rect 12256 12106 12308 12112
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12452 11354 12480 11766
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9926 12480 10066
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 12544 9586 12572 12582
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12636 11558 12664 12378
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12636 10062 12664 11494
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12728 9586 12756 12038
rect 12820 11694 12848 12718
rect 12912 12442 12940 13330
rect 13004 12918 13032 13330
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 13004 11218 13032 12718
rect 13096 11830 13124 13330
rect 13188 12442 13216 13330
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12918 13860 13126
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 14108 12850 14136 13466
rect 14476 13394 14504 13806
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 15028 13394 15056 13942
rect 15212 13802 15240 14350
rect 15304 14006 15332 14418
rect 15764 14414 15792 16594
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15856 14482 15884 14826
rect 16592 14550 16620 15846
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 16900 15260 17208 15269
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 17512 15026 17540 15438
rect 18340 15094 18368 15438
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 16960 14414 16988 14962
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15304 13394 15332 13942
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 13394 15608 13738
rect 16224 13462 16252 13806
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 12850 14320 13194
rect 14556 13184 14608 13190
rect 14476 13144 14556 13172
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13556 12594 13584 12650
rect 13372 12566 13584 12594
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13372 12238 13400 12566
rect 14476 12434 14504 13144
rect 14556 13126 14608 13132
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 14384 12406 14504 12434
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 12102 13400 12174
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 13372 11558 13400 12038
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 11286 13400 11494
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12820 11121 12848 11154
rect 12806 11112 12862 11121
rect 12806 11047 12862 11056
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12820 9586 12848 10066
rect 12992 10056 13044 10062
rect 12898 10024 12954 10033
rect 12992 9998 13044 10004
rect 12898 9959 12954 9968
rect 12912 9586 12940 9959
rect 13004 9722 13032 9998
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12176 8906 12204 9046
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12544 8537 12572 9318
rect 12820 9178 12848 9318
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12716 8968 12768 8974
rect 12912 8945 12940 9386
rect 12716 8910 12768 8916
rect 12898 8936 12954 8945
rect 12530 8528 12586 8537
rect 11900 8486 12204 8514
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11624 6866 11652 6938
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11716 6662 11744 7142
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11426 5879 11482 5888
rect 11520 5908 11572 5914
rect 11440 5846 11468 5879
rect 11520 5850 11572 5856
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 3670 11376 4966
rect 11440 4826 11468 5782
rect 11624 5302 11652 6598
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11532 4146 11560 4966
rect 11624 4690 11652 5238
rect 11716 4826 11744 6598
rect 11808 5794 11836 6870
rect 11900 6730 11928 8366
rect 12176 8362 12204 8486
rect 12530 8463 12586 8472
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12452 8294 12480 8366
rect 12440 8288 12492 8294
rect 12162 8256 12218 8265
rect 12440 8230 12492 8236
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12162 8191 12218 8200
rect 12176 7954 12204 8191
rect 12452 7993 12480 8230
rect 12438 7984 12494 7993
rect 12164 7948 12216 7954
rect 12438 7919 12440 7928
rect 12164 7890 12216 7896
rect 12492 7919 12494 7928
rect 12440 7890 12492 7896
rect 12438 7848 12494 7857
rect 12438 7783 12440 7792
rect 12492 7783 12494 7792
rect 12440 7754 12492 7760
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11808 5766 11928 5794
rect 11992 5778 12020 7686
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 12544 7478 12572 8230
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11808 4826 11836 5646
rect 11900 5352 11928 5766
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11900 5324 12020 5352
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 10980 2746 11284 2774
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10416 1556 10468 1562
rect 10416 1498 10468 1504
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 10704 1358 10732 2382
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 10888 1358 10916 1838
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 10876 1352 10928 1358
rect 10876 1294 10928 1300
rect 10888 882 10916 1294
rect 10876 876 10928 882
rect 10876 818 10928 824
rect 9404 808 9456 814
rect 9404 750 9456 756
rect 8668 740 8720 746
rect 8668 682 8720 688
rect 7288 672 7340 678
rect 7288 614 7340 620
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 3896 462 4016 490
rect 3896 400 3924 462
rect 10980 400 11008 2746
rect 11440 2428 11468 2994
rect 11532 2990 11560 3878
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11716 2922 11744 4014
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11612 2440 11664 2446
rect 11440 2400 11612 2428
rect 11612 2382 11664 2388
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 1426 11560 2246
rect 11624 1970 11652 2382
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 11716 1766 11744 2858
rect 11808 2106 11836 4762
rect 11900 4128 11928 5170
rect 11992 5166 12020 5324
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11992 5030 12020 5102
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11980 4140 12032 4146
rect 11900 4100 11980 4128
rect 11980 4082 12032 4088
rect 11992 3058 12020 4082
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11992 1902 12020 2382
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11992 1494 12020 1702
rect 11980 1488 12032 1494
rect 11980 1430 12032 1436
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11992 814 12020 1430
rect 12084 898 12112 7210
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12360 6662 12388 6802
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 12544 6186 12572 6802
rect 12636 6390 12664 7754
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 5681 12388 5714
rect 12346 5672 12402 5681
rect 12346 5607 12402 5616
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 12544 5370 12572 6122
rect 12728 5778 12756 8910
rect 12898 8871 12954 8880
rect 13280 8838 13308 9862
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12992 8424 13044 8430
rect 12820 8384 12992 8412
rect 12820 6730 12848 8384
rect 12992 8366 13044 8372
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 8129 13032 8230
rect 12990 8120 13046 8129
rect 12990 8055 13046 8064
rect 13004 7954 13032 8055
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12900 7880 12952 7886
rect 12898 7848 12900 7857
rect 12952 7848 12954 7857
rect 13188 7834 13216 7890
rect 12954 7806 13216 7834
rect 12898 7783 12954 7792
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7206 13124 7686
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12806 6624 12862 6633
rect 12806 6559 12862 6568
rect 12820 6186 12848 6559
rect 12912 6254 12940 6802
rect 13188 6662 13216 7806
rect 13372 7478 13400 8978
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13174 6352 13230 6361
rect 13174 6287 13176 6296
rect 13228 6287 13230 6296
rect 13176 6258 13228 6264
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12716 5772 12768 5778
rect 12636 5732 12716 5760
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12268 4826 12296 5102
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12176 4486 12204 4694
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 12544 3534 12572 4558
rect 12636 4214 12664 5732
rect 12716 5714 12768 5720
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5234 12756 5510
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12820 4282 12848 6122
rect 12992 6112 13044 6118
rect 12990 6080 12992 6089
rect 13044 6080 13046 6089
rect 12990 6015 13046 6024
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5166 13032 5510
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 13004 3534 13032 4966
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 13280 2774 13308 7210
rect 13372 6254 13400 7414
rect 13464 6730 13492 7686
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13556 6254 13584 11630
rect 13832 11286 13860 12310
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13832 10538 13860 11018
rect 13924 10742 13952 11018
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13832 10266 13860 10474
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13832 10130 13860 10202
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13924 9994 13952 10678
rect 14016 10606 14044 12174
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11218 14228 11494
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14200 10538 14228 11154
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14200 10266 14228 10474
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14108 9042 14136 9590
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13726 7984 13782 7993
rect 13636 7948 13688 7954
rect 13782 7928 13860 7936
rect 13726 7919 13728 7928
rect 13636 7890 13688 7896
rect 13780 7908 13860 7928
rect 13728 7890 13780 7896
rect 13648 7818 13676 7890
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13648 7177 13676 7754
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13740 7313 13768 7414
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 13634 7168 13690 7177
rect 13634 7103 13690 7112
rect 13832 6934 13860 7908
rect 13924 7449 13952 8366
rect 14016 7818 14044 8434
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13910 7440 13966 7449
rect 13910 7375 13966 7384
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13726 6760 13782 6769
rect 13648 6718 13726 6746
rect 13360 6248 13412 6254
rect 13358 6216 13360 6225
rect 13544 6248 13596 6254
rect 13412 6216 13414 6225
rect 13544 6190 13596 6196
rect 13358 6151 13414 6160
rect 13648 6089 13676 6718
rect 13726 6695 13782 6704
rect 13832 6458 13860 6870
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13634 6080 13690 6089
rect 13634 6015 13690 6024
rect 13648 5778 13676 6015
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13372 5370 13400 5646
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 5030 13400 5306
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13740 4622 13768 5510
rect 13832 5302 13860 6122
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13740 3738 13768 4014
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13924 2854 13952 7375
rect 14108 7342 14136 7482
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14002 7168 14058 7177
rect 14002 7103 14058 7112
rect 14016 6798 14044 7103
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14200 6458 14228 10066
rect 14384 9518 14412 12406
rect 15120 12306 15148 12718
rect 15304 12646 15332 13330
rect 15580 12918 15608 13330
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15120 12170 15148 12242
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 11762 15148 12106
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15106 11656 15162 11665
rect 15106 11591 15108 11600
rect 15160 11591 15162 11600
rect 15108 11562 15160 11568
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 15028 11150 15056 11494
rect 15212 11218 15240 12378
rect 15580 12306 15608 12854
rect 16224 12850 16252 13398
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 16500 12238 16528 12718
rect 16684 12442 16712 14214
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 15304 11694 15332 12174
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10713 14780 10950
rect 14738 10704 14794 10713
rect 14738 10639 14794 10648
rect 14844 10606 14872 11018
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14936 10606 14964 10678
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14542 10299 14850 10308
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14476 9722 14504 9998
rect 14936 9926 14964 10542
rect 15028 10130 15056 10610
rect 15212 10606 15240 11154
rect 15304 10674 15332 11222
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15108 10464 15160 10470
rect 15580 10418 15608 10610
rect 16316 10606 16344 12038
rect 16500 11694 16528 12174
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 17328 11694 17356 14418
rect 17512 13530 17540 14962
rect 18340 14482 18368 15030
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18340 14346 18368 14418
rect 18880 14408 18932 14414
rect 18984 14385 19012 16594
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19076 15065 19104 15982
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 19062 15056 19118 15065
rect 19062 14991 19118 15000
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 18880 14350 18932 14356
rect 18970 14376 19026 14385
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 17604 13870 17632 14282
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17604 13394 17632 13806
rect 18708 13734 18736 14214
rect 18892 14074 18920 14350
rect 18970 14311 19026 14320
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17880 12646 17908 13194
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12306 17908 12582
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17880 12170 17908 12242
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11694 17908 12106
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 16500 11218 16528 11630
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10674 16528 11154
rect 17144 11014 17172 11562
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 16488 10668 16540 10674
rect 16540 10628 16620 10656
rect 16488 10610 16540 10616
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 15108 10406 15160 10412
rect 15120 10146 15148 10406
rect 15212 10390 15608 10418
rect 15212 10266 15240 10390
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15120 10130 15240 10146
rect 15016 10124 15068 10130
rect 15120 10124 15252 10130
rect 15120 10118 15200 10124
rect 15016 10066 15068 10072
rect 15396 10112 15424 10202
rect 15580 10130 15608 10390
rect 15948 10266 15976 10474
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15568 10124 15620 10130
rect 15396 10084 15516 10112
rect 15200 10066 15252 10072
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14660 9518 14688 9862
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14476 9178 14504 9454
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14292 8430 14320 8978
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8430 14504 8910
rect 14936 8650 14964 9318
rect 15028 9042 15056 9930
rect 15120 9518 15148 9998
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15488 9976 15516 10084
rect 15568 10066 15620 10072
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15568 9988 15620 9994
rect 15488 9948 15568 9976
rect 15212 9874 15240 9930
rect 15290 9888 15346 9897
rect 15212 9846 15290 9874
rect 15290 9823 15346 9832
rect 15488 9602 15516 9948
rect 15568 9930 15620 9936
rect 15672 9722 15700 10066
rect 15750 10024 15806 10033
rect 15750 9959 15806 9968
rect 16120 9988 16172 9994
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15304 9574 15516 9602
rect 15566 9616 15622 9625
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 9042 15148 9454
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14752 8622 14964 8650
rect 14752 8498 14780 8622
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14292 6633 14320 7278
rect 14384 6934 14412 7754
rect 14568 7478 14596 7754
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14094 6216 14150 6225
rect 14094 6151 14150 6160
rect 14108 5778 14136 6151
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14108 5302 14136 5714
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14016 4146 14044 5034
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13188 2746 13308 2774
rect 13188 2514 13216 2746
rect 14108 2514 14136 2926
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 12636 1358 12664 2450
rect 14108 1970 14136 2450
rect 14200 2038 14228 6394
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14292 5030 14320 6258
rect 14384 6254 14412 6870
rect 14936 6769 14964 8622
rect 15212 8430 15240 9522
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 15028 7954 15056 8298
rect 15120 7954 15148 8366
rect 15304 8294 15332 9574
rect 15764 9586 15792 9959
rect 16120 9930 16172 9936
rect 15844 9920 15896 9926
rect 15842 9888 15844 9897
rect 15896 9888 15898 9897
rect 15842 9823 15898 9832
rect 15566 9551 15622 9560
rect 15752 9580 15804 9586
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 8498 15424 9454
rect 15580 9110 15608 9551
rect 15752 9522 15804 9528
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 14922 6760 14978 6769
rect 14922 6695 14978 6704
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14476 2922 14504 6190
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 15028 5658 15056 7754
rect 15120 6798 15148 7890
rect 15200 6928 15252 6934
rect 15198 6896 15200 6905
rect 15252 6896 15254 6905
rect 15304 6866 15332 8230
rect 15396 7410 15424 8434
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15198 6831 15254 6840
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15396 6730 15424 7346
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15488 5914 15516 6734
rect 15580 5914 15608 6938
rect 15672 6458 15700 8978
rect 16132 8838 16160 9930
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16224 8430 16252 10474
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10130 16528 10406
rect 16592 10130 16620 10628
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9518 16436 9862
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16408 9110 16436 9454
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16500 8906 16528 10066
rect 16776 9042 16804 10066
rect 16900 9820 17208 9829
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 17236 9042 17264 10066
rect 17328 10062 17356 11494
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17420 10985 17448 11290
rect 17880 11082 17908 11630
rect 18248 11286 18276 13330
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12850 18644 13126
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18892 12238 18920 13806
rect 18984 12322 19012 14214
rect 19076 14113 19104 14826
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 19062 14104 19118 14113
rect 19062 14039 19118 14048
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19168 13025 19196 13806
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 19154 13016 19210 13025
rect 19154 12951 19210 12960
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 19062 12336 19118 12345
rect 18984 12294 19062 12322
rect 19062 12271 19118 12280
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11286 18920 12174
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17406 10976 17462 10985
rect 17406 10911 17462 10920
rect 17880 10674 17908 11018
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16408 7954 16436 8366
rect 16592 7954 16620 8502
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15856 6866 15884 7278
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15672 6361 15700 6394
rect 15658 6352 15714 6361
rect 15764 6322 15792 6666
rect 15658 6287 15714 6296
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 6186 15792 6258
rect 15856 6254 15884 6802
rect 15948 6662 15976 7890
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16670 7304 16726 7313
rect 16040 6730 16068 7278
rect 16670 7239 16726 7248
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16040 6322 16068 6666
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15106 5672 15162 5681
rect 15028 5630 15106 5658
rect 15290 5672 15346 5681
rect 15106 5607 15162 5616
rect 15212 5630 15290 5658
rect 15212 5574 15240 5630
rect 15290 5607 15346 5616
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15292 5568 15344 5574
rect 15396 5545 15424 5714
rect 15764 5642 15792 6122
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15292 5510 15344 5516
rect 15382 5536 15438 5545
rect 15304 5166 15332 5510
rect 15382 5471 15438 5480
rect 15396 5166 15424 5471
rect 15764 5302 15792 5578
rect 15856 5302 15884 5714
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 15396 4690 15424 5102
rect 15672 5098 15700 5238
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15948 4690 15976 5714
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14844 4214 14872 4490
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 14936 3670 14964 4422
rect 16040 4196 16068 6258
rect 16302 5808 16358 5817
rect 16408 5778 16436 6666
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16302 5743 16358 5752
rect 16396 5772 16448 5778
rect 16316 5710 16344 5743
rect 16396 5714 16448 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16132 5370 16160 5510
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16132 4826 16160 5306
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16224 4826 16252 5238
rect 16316 5166 16344 5646
rect 16408 5545 16436 5714
rect 16394 5536 16450 5545
rect 16394 5471 16450 5480
rect 16592 5166 16620 6598
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 15474 4176 15530 4185
rect 16040 4168 16252 4196
rect 15474 4111 15530 4120
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 14542 2683 14850 2692
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14188 2032 14240 2038
rect 14188 1974 14240 1980
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 13648 1426 13676 1906
rect 14476 1902 14504 2314
rect 14464 1896 14516 1902
rect 14464 1838 14516 1844
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 13636 1420 13688 1426
rect 13636 1362 13688 1368
rect 12624 1352 12676 1358
rect 12624 1294 12676 1300
rect 13452 1352 13504 1358
rect 13452 1294 13504 1300
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 12084 870 12296 898
rect 13464 882 13492 1294
rect 13648 950 13676 1362
rect 13636 944 13688 950
rect 13636 886 13688 892
rect 14936 882 14964 3062
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 15028 1902 15056 2042
rect 15016 1896 15068 1902
rect 15016 1838 15068 1844
rect 11980 808 12032 814
rect 11980 750 12032 756
rect 12268 400 12296 870
rect 13452 876 13504 882
rect 13452 818 13504 824
rect 14924 876 14976 882
rect 14924 818 14976 824
rect 15028 814 15056 1838
rect 15488 1426 15516 4111
rect 16224 4010 16252 4168
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16224 3194 16252 3946
rect 16316 3738 16344 4626
rect 16500 4622 16528 5034
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15764 1494 15792 2382
rect 15856 1902 15884 2450
rect 16224 2038 16252 2994
rect 16592 2650 16620 5102
rect 16684 4758 16712 7239
rect 16776 6934 16804 8978
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16854 6896 16910 6905
rect 16854 6831 16856 6840
rect 16908 6831 16910 6840
rect 16856 6802 16908 6808
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16776 6322 16804 6666
rect 16868 6662 16896 6802
rect 17236 6662 17264 8978
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16684 4078 16712 4150
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16776 3194 16804 6258
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16960 5642 16988 6122
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5778 17264 6054
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 17328 5114 17356 9998
rect 17420 8498 17448 10406
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 8974 17540 10066
rect 17972 10062 18000 10542
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17604 8430 17632 9454
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17604 7954 17632 8366
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17696 7342 17724 9454
rect 17880 9042 17908 9454
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17788 7818 17816 8434
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7410 17816 7754
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17406 6760 17462 6769
rect 17406 6695 17462 6704
rect 17144 5086 17356 5114
rect 17420 5098 17448 6695
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17512 6322 17540 6394
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17604 6186 17632 6870
rect 17592 6180 17644 6186
rect 17592 6122 17644 6128
rect 17696 5914 17724 7278
rect 17788 6798 17816 7346
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17408 5092 17460 5098
rect 17144 4690 17172 5086
rect 17408 5034 17460 5040
rect 17224 5024 17276 5030
rect 17420 4978 17448 5034
rect 17224 4966 17276 4972
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 17236 4078 17264 4966
rect 17328 4950 17448 4978
rect 17328 4690 17356 4950
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16212 2032 16264 2038
rect 16212 1974 16264 1980
rect 16776 1970 16804 3130
rect 17236 3058 17264 4014
rect 17420 3602 17448 4762
rect 17512 3738 17540 5102
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17604 3602 17632 5102
rect 17788 4282 17816 6190
rect 17880 4826 17908 8298
rect 18064 7478 18092 9590
rect 18156 9586 18184 10406
rect 18248 9722 18276 11222
rect 19076 11054 19104 11630
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 19076 11026 19196 11054
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 7478 18184 9318
rect 18432 8974 18460 9998
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18524 9586 18552 9930
rect 18708 9722 18736 10542
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18248 7954 18276 8230
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18340 7478 18368 8570
rect 18432 8566 18460 8910
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18616 8090 18644 8842
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6254 18000 6598
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 18064 5710 18092 7414
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18064 5098 18092 5646
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 18064 4214 18092 4558
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 18064 3210 18092 4150
rect 18156 3602 18184 6802
rect 18248 6458 18276 7210
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 17926 3182 18092 3210
rect 17926 3108 17954 3182
rect 17880 3080 17954 3108
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 16764 1964 16816 1970
rect 16764 1906 16816 1912
rect 15844 1896 15896 1902
rect 15844 1838 15896 1844
rect 15752 1488 15804 1494
rect 15752 1430 15804 1436
rect 17512 1426 17540 2858
rect 17880 2378 17908 3080
rect 18064 3058 18092 3182
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 17880 2038 17908 2314
rect 17868 2032 17920 2038
rect 17868 1974 17920 1980
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 17500 1420 17552 1426
rect 17500 1362 17552 1368
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16132 882 16160 1294
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 16120 876 16172 882
rect 16120 818 16172 824
rect 17512 814 17540 1362
rect 17880 1358 17908 1974
rect 17972 1902 18000 2926
rect 18340 2514 18368 6258
rect 18432 6254 18460 8026
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 5370 18460 6054
rect 18524 5778 18552 7890
rect 18708 7546 18736 8230
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18616 6390 18644 6802
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18616 5846 18644 6326
rect 18708 6322 18736 7142
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18800 6254 18828 9386
rect 18892 8566 18920 9454
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18892 7546 18920 8502
rect 18984 7954 19012 9862
rect 19076 8945 19104 10406
rect 19062 8936 19118 8945
rect 19062 8871 19118 8880
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18788 6248 18840 6254
rect 18694 6216 18750 6225
rect 18788 6190 18840 6196
rect 18694 6151 18750 6160
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18524 5166 18552 5578
rect 18602 5536 18658 5545
rect 18602 5471 18658 5480
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4622 18552 5102
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18616 3602 18644 5471
rect 18708 4078 18736 6151
rect 18892 5778 18920 7278
rect 18984 6202 19012 7890
rect 19062 7576 19118 7585
rect 19168 7562 19196 11026
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 19706 7848 19762 7857
rect 19706 7783 19762 7792
rect 19118 7534 19196 7562
rect 19062 7511 19118 7520
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 19430 6896 19486 6905
rect 19486 6854 19656 6882
rect 19430 6831 19486 6840
rect 18984 6174 19196 6202
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18972 5704 19024 5710
rect 18786 5672 18842 5681
rect 18972 5646 19024 5652
rect 18786 5607 18842 5616
rect 18800 5166 18828 5607
rect 18984 5166 19012 5646
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 19076 4154 19104 6054
rect 19168 4690 19196 6174
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18892 4126 19104 4154
rect 18892 4078 18920 4126
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 19628 2514 19656 6854
rect 19720 2990 19748 7783
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 19614 2408 19670 2417
rect 17960 1896 18012 1902
rect 17960 1838 18012 1844
rect 18248 1426 18276 2382
rect 19614 2343 19670 2352
rect 19062 2136 19118 2145
rect 19062 2071 19118 2080
rect 18880 1896 18932 1902
rect 18880 1838 18932 1844
rect 18512 1760 18564 1766
rect 18512 1702 18564 1708
rect 18524 1494 18552 1702
rect 18512 1488 18564 1494
rect 18892 1465 18920 1838
rect 18512 1430 18564 1436
rect 18878 1456 18934 1465
rect 18236 1420 18288 1426
rect 18878 1391 18934 1400
rect 18236 1362 18288 1368
rect 17868 1352 17920 1358
rect 17868 1294 17920 1300
rect 17880 950 17908 1294
rect 19076 1018 19104 2071
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 19628 1426 19656 2343
rect 19616 1420 19668 1426
rect 19616 1362 19668 1368
rect 19064 1012 19116 1018
rect 19064 954 19116 960
rect 17868 944 17920 950
rect 17868 886 17920 892
rect 15016 808 15068 814
rect 15016 750 15068 756
rect 17500 808 17552 814
rect 17500 750 17552 756
rect 15476 672 15528 678
rect 15476 614 15528 620
rect 18052 672 18104 678
rect 18052 614 18104 620
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 15488 400 15516 614
rect 18064 400 18092 614
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 18 0 74 400
rect 662 0 718 400
rect 1306 0 1362 400
rect 1950 0 2006 400
rect 2594 0 2650 400
rect 3882 0 3938 400
rect 10966 0 11022 400
rect 12254 0 12310 400
rect 15474 0 15530 400
rect 18050 0 18106 400
<< via2 >>
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 846 18400 902 18456
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 3606 17720 3662 17776
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 4342 6296 4398 6352
rect 4618 6160 4674 6216
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 478 4120 534 4176
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 5170 6316 5226 6352
rect 5170 6296 5172 6316
rect 5172 6296 5224 6316
rect 5224 6296 5226 6316
rect 5446 6160 5502 6216
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 8298 13096 8354 13152
rect 8022 12300 8078 12336
rect 8022 12280 8024 12300
rect 8024 12280 8076 12300
rect 8076 12280 8078 12300
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 7838 8880 7894 8936
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 8390 10668 8446 10704
rect 8390 10648 8392 10668
rect 8392 10648 8444 10668
rect 8444 10648 8446 10668
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 8942 13368 8998 13424
rect 8942 13252 8998 13288
rect 8942 13232 8944 13252
rect 8944 13232 8996 13252
rect 8996 13232 8998 13252
rect 8758 12688 8814 12744
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 9586 15272 9642 15328
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 9126 12316 9128 12336
rect 9128 12316 9180 12336
rect 9180 12316 9182 12336
rect 9126 12280 9182 12316
rect 9126 10920 9182 10976
rect 9862 13252 9918 13288
rect 9862 13232 9864 13252
rect 9864 13232 9916 13252
rect 9916 13232 9918 13252
rect 10230 12688 10286 12744
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 10046 11600 10102 11656
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 10046 11212 10102 11248
rect 10046 11192 10048 11212
rect 10048 11192 10100 11212
rect 10100 11192 10102 11212
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 10046 10668 10102 10704
rect 10046 10648 10048 10668
rect 10048 10648 10100 10668
rect 10100 10648 10102 10668
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 10782 12844 10838 12880
rect 10782 12824 10784 12844
rect 10784 12824 10836 12844
rect 10836 12824 10838 12844
rect 10690 12144 10746 12200
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 9770 9832 9826 9888
rect 10138 9988 10194 10024
rect 10138 9968 10140 9988
rect 10140 9968 10192 9988
rect 10192 9968 10194 9988
rect 10046 9832 10102 9888
rect 10230 9696 10286 9752
rect 10138 9460 10140 9480
rect 10140 9460 10192 9480
rect 10192 9460 10194 9480
rect 10138 9424 10194 9460
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 9862 8880 9918 8936
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 10506 8880 10562 8936
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 8482 4120 8538 4176
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 846 1400 902 1456
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 11058 12316 11060 12336
rect 11060 12316 11112 12336
rect 11112 12316 11114 12336
rect 11058 12280 11114 12316
rect 11058 9696 11114 9752
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 11426 13096 11482 13152
rect 11610 12280 11666 12336
rect 11426 9696 11482 9752
rect 10966 9424 11022 9480
rect 11150 9424 11206 9480
rect 11150 8472 11206 8528
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 11518 8064 11574 8120
rect 11426 5888 11482 5944
rect 11702 8200 11758 8256
rect 11702 7384 11758 7440
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 12162 13388 12218 13424
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 12162 13368 12164 13388
rect 12164 13368 12216 13388
rect 12216 13368 12218 13388
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 12254 12280 12310 12336
rect 12346 12144 12402 12200
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 12806 11056 12862 11112
rect 12898 9968 12954 10024
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 12530 8472 12586 8528
rect 12162 8200 12218 8256
rect 12438 7948 12494 7984
rect 12438 7928 12440 7948
rect 12440 7928 12492 7948
rect 12492 7928 12494 7948
rect 12438 7812 12494 7848
rect 12438 7792 12440 7812
rect 12440 7792 12492 7812
rect 12492 7792 12494 7812
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 12346 5616 12402 5672
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 12898 8880 12954 8936
rect 12990 8064 13046 8120
rect 12898 7828 12900 7848
rect 12900 7828 12952 7848
rect 12952 7828 12954 7848
rect 12898 7792 12954 7828
rect 12806 6568 12862 6624
rect 13174 6316 13230 6352
rect 13174 6296 13176 6316
rect 13176 6296 13228 6316
rect 13228 6296 13230 6316
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 12990 6060 12992 6080
rect 12992 6060 13044 6080
rect 13044 6060 13046 6080
rect 12990 6024 13046 6060
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 13726 7948 13782 7984
rect 13726 7928 13728 7948
rect 13728 7928 13780 7948
rect 13780 7928 13782 7948
rect 13726 7248 13782 7304
rect 13634 7112 13690 7168
rect 13910 7384 13966 7440
rect 13358 6196 13360 6216
rect 13360 6196 13412 6216
rect 13412 6196 13414 6216
rect 13358 6160 13414 6196
rect 13726 6704 13782 6760
rect 13634 6024 13690 6080
rect 14002 7112 14058 7168
rect 15106 11620 15162 11656
rect 15106 11600 15108 11620
rect 15108 11600 15160 11620
rect 15160 11600 15162 11620
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 14738 10648 14794 10704
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 19062 15000 19118 15056
rect 18970 14320 19026 14376
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 15290 9832 15346 9888
rect 15750 9968 15806 10024
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 14278 6568 14334 6624
rect 14094 6160 14150 6216
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 15566 9560 15622 9616
rect 15842 9868 15844 9888
rect 15844 9868 15896 9888
rect 15896 9868 15898 9888
rect 15842 9832 15898 9868
rect 14922 6704 14978 6760
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 15198 6876 15200 6896
rect 15200 6876 15252 6896
rect 15252 6876 15254 6896
rect 15198 6840 15254 6876
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 19062 14048 19118 14104
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 19154 12960 19210 13016
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 19062 12280 19118 12336
rect 17406 10920 17462 10976
rect 15658 6296 15714 6352
rect 16670 7248 16726 7304
rect 15106 5616 15162 5672
rect 15290 5616 15346 5672
rect 15382 5480 15438 5536
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 16302 5752 16358 5808
rect 16394 5480 16450 5536
rect 15474 4120 15530 4176
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 16854 6860 16910 6896
rect 16854 6840 16856 6860
rect 16856 6840 16908 6860
rect 16908 6840 16910 6860
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 17406 6704 17462 6760
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 19062 8880 19118 8936
rect 18694 6160 18750 6216
rect 18602 5480 18658 5536
rect 19062 7520 19118 7576
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 19706 7792 19762 7848
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 19430 6840 19486 6896
rect 18786 5616 18842 5672
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 19614 2352 19670 2408
rect 19062 2080 19118 2136
rect 18878 1400 18934 1456
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
<< metal3 >>
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19253 19007 19569 19008
rect 2751 18528 3067 18529
rect 0 18458 400 18488
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 841 18458 907 18461
rect 0 18456 907 18458
rect 0 18400 846 18456
rect 902 18400 907 18456
rect 0 18398 907 18400
rect 0 18368 400 18398
rect 841 18395 907 18398
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 0 17778 400 17808
rect 3601 17778 3667 17781
rect 0 17776 3667 17778
rect 0 17720 3606 17776
rect 3662 17720 3667 17776
rect 0 17718 3667 17720
rect 0 17688 400 17718
rect 3601 17715 3667 17718
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 9254 15268 9260 15332
rect 9324 15330 9330 15332
rect 9581 15330 9647 15333
rect 9324 15328 9647 15330
rect 9324 15272 9586 15328
rect 9642 15272 9647 15328
rect 9324 15270 9647 15272
rect 9324 15268 9330 15270
rect 9581 15267 9647 15270
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 19057 15058 19123 15061
rect 19600 15058 20000 15088
rect 19057 15056 20000 15058
rect 19057 15000 19062 15056
rect 19118 15000 20000 15056
rect 19057 14998 20000 15000
rect 19057 14995 19123 14998
rect 19600 14968 20000 14998
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 18965 14378 19031 14381
rect 19600 14378 20000 14408
rect 18965 14376 20000 14378
rect 18965 14320 18970 14376
rect 19026 14320 20000 14376
rect 18965 14318 20000 14320
rect 18965 14315 19031 14318
rect 19600 14288 20000 14318
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 19057 14106 19123 14109
rect 19057 14104 19810 14106
rect 19057 14048 19062 14104
rect 19118 14048 19810 14104
rect 19057 14046 19810 14048
rect 19057 14043 19123 14046
rect 19750 13728 19810 14046
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19600 13608 20000 13728
rect 19253 13567 19569 13568
rect 8937 13426 9003 13429
rect 12157 13426 12223 13429
rect 8937 13424 12223 13426
rect 8937 13368 8942 13424
rect 8998 13368 12162 13424
rect 12218 13368 12223 13424
rect 8937 13366 12223 13368
rect 8937 13363 9003 13366
rect 12157 13363 12223 13366
rect 8937 13290 9003 13293
rect 9857 13290 9923 13293
rect 8937 13288 9923 13290
rect 8937 13232 8942 13288
rect 8998 13232 9862 13288
rect 9918 13232 9923 13288
rect 8937 13230 9923 13232
rect 8937 13227 9003 13230
rect 9857 13227 9923 13230
rect 8293 13154 8359 13157
rect 11421 13154 11487 13157
rect 8293 13152 11487 13154
rect 8293 13096 8298 13152
rect 8354 13096 11426 13152
rect 11482 13096 11487 13152
rect 8293 13094 11487 13096
rect 8293 13091 8359 13094
rect 11421 13091 11487 13094
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 19149 13018 19215 13021
rect 19600 13018 20000 13048
rect 19149 13016 20000 13018
rect 19149 12960 19154 13016
rect 19210 12960 20000 13016
rect 19149 12958 20000 12960
rect 19149 12955 19215 12958
rect 19600 12928 20000 12958
rect 9622 12820 9628 12884
rect 9692 12882 9698 12884
rect 10777 12882 10843 12885
rect 9692 12880 10843 12882
rect 9692 12824 10782 12880
rect 10838 12824 10843 12880
rect 9692 12822 10843 12824
rect 9692 12820 9698 12822
rect 10777 12819 10843 12822
rect 8753 12746 8819 12749
rect 10225 12746 10291 12749
rect 8753 12744 10291 12746
rect 8753 12688 8758 12744
rect 8814 12688 10230 12744
rect 10286 12688 10291 12744
rect 8753 12686 10291 12688
rect 8753 12683 8819 12686
rect 10225 12683 10291 12686
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 8017 12338 8083 12341
rect 9121 12338 9187 12341
rect 8017 12336 9187 12338
rect 8017 12280 8022 12336
rect 8078 12280 9126 12336
rect 9182 12280 9187 12336
rect 8017 12278 9187 12280
rect 8017 12275 8083 12278
rect 9121 12275 9187 12278
rect 11053 12338 11119 12341
rect 11605 12338 11671 12341
rect 12249 12338 12315 12341
rect 11053 12336 12315 12338
rect 11053 12280 11058 12336
rect 11114 12280 11610 12336
rect 11666 12280 12254 12336
rect 12310 12280 12315 12336
rect 11053 12278 12315 12280
rect 11053 12275 11119 12278
rect 11605 12275 11671 12278
rect 12249 12275 12315 12278
rect 19057 12338 19123 12341
rect 19600 12338 20000 12368
rect 19057 12336 20000 12338
rect 19057 12280 19062 12336
rect 19118 12280 20000 12336
rect 19057 12278 20000 12280
rect 19057 12275 19123 12278
rect 19600 12248 20000 12278
rect 10685 12202 10751 12205
rect 12341 12202 12407 12205
rect 10685 12200 12407 12202
rect 10685 12144 10690 12200
rect 10746 12144 12346 12200
rect 12402 12144 12407 12200
rect 10685 12142 12407 12144
rect 10685 12139 10751 12142
rect 12341 12139 12407 12142
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 10041 11658 10107 11661
rect 15101 11658 15167 11661
rect 19600 11658 20000 11688
rect 10041 11656 10288 11658
rect 10041 11600 10046 11656
rect 10102 11600 10288 11656
rect 10041 11598 10288 11600
rect 10041 11595 10107 11598
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 10041 11250 10107 11253
rect 10228 11250 10288 11598
rect 15101 11656 20000 11658
rect 15101 11600 15106 11656
rect 15162 11600 20000 11656
rect 15101 11598 20000 11600
rect 15101 11595 15167 11598
rect 19600 11568 20000 11598
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 10041 11248 10288 11250
rect 10041 11192 10046 11248
rect 10102 11192 10288 11248
rect 10041 11190 10288 11192
rect 10041 11187 10107 11190
rect 12566 11052 12572 11116
rect 12636 11114 12642 11116
rect 12801 11114 12867 11117
rect 12636 11112 12867 11114
rect 12636 11056 12806 11112
rect 12862 11056 12867 11112
rect 12636 11054 12867 11056
rect 12636 11052 12642 11054
rect 12801 11051 12867 11054
rect 0 10978 400 11008
rect 9121 10978 9187 10981
rect 9254 10978 9260 10980
rect 0 10918 1410 10978
rect 0 10888 400 10918
rect 1350 10706 1410 10918
rect 9121 10976 9260 10978
rect 9121 10920 9126 10976
rect 9182 10920 9260 10976
rect 9121 10918 9260 10920
rect 9121 10915 9187 10918
rect 9254 10916 9260 10918
rect 9324 10916 9330 10980
rect 17401 10978 17467 10981
rect 19600 10978 20000 11008
rect 17401 10976 20000 10978
rect 17401 10920 17406 10976
rect 17462 10920 20000 10976
rect 17401 10918 20000 10920
rect 17401 10915 17467 10918
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 19600 10888 20000 10918
rect 16896 10847 17212 10848
rect 8385 10706 8451 10709
rect 1350 10704 8451 10706
rect 1350 10648 8390 10704
rect 8446 10648 8451 10704
rect 1350 10646 8451 10648
rect 8385 10643 8451 10646
rect 10041 10706 10107 10709
rect 14733 10706 14799 10709
rect 10041 10704 14799 10706
rect 10041 10648 10046 10704
rect 10102 10648 14738 10704
rect 14794 10648 14799 10704
rect 10041 10646 14799 10648
rect 10041 10643 10107 10646
rect 14733 10643 14799 10646
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 19600 10208 20000 10328
rect 10133 10026 10199 10029
rect 12893 10026 12959 10029
rect 10133 10024 12959 10026
rect 10133 9968 10138 10024
rect 10194 9968 12898 10024
rect 12954 9968 12959 10024
rect 10133 9966 12959 9968
rect 10133 9963 10199 9966
rect 12893 9963 12959 9966
rect 15745 10026 15811 10029
rect 19750 10026 19810 10208
rect 15745 10024 19810 10026
rect 15745 9968 15750 10024
rect 15806 9968 19810 10024
rect 15745 9966 19810 9968
rect 15745 9963 15811 9966
rect 9765 9890 9831 9893
rect 10041 9890 10107 9893
rect 9765 9888 10107 9890
rect 9765 9832 9770 9888
rect 9826 9832 10046 9888
rect 10102 9832 10107 9888
rect 9765 9830 10107 9832
rect 9765 9827 9831 9830
rect 10041 9827 10107 9830
rect 15285 9890 15351 9893
rect 15837 9890 15903 9893
rect 15285 9888 15903 9890
rect 15285 9832 15290 9888
rect 15346 9832 15842 9888
rect 15898 9832 15903 9888
rect 15285 9830 15903 9832
rect 15285 9827 15351 9830
rect 15837 9827 15903 9830
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 16896 9759 17212 9760
rect 10225 9754 10291 9757
rect 11053 9754 11119 9757
rect 11421 9754 11487 9757
rect 10225 9752 11119 9754
rect 10225 9696 10230 9752
rect 10286 9696 11058 9752
rect 11114 9696 11119 9752
rect 10225 9694 11119 9696
rect 10225 9691 10291 9694
rect 11053 9691 11119 9694
rect 11286 9752 11487 9754
rect 11286 9696 11426 9752
rect 11482 9696 11487 9752
rect 11286 9694 11487 9696
rect 10133 9482 10199 9485
rect 10961 9482 11027 9485
rect 10133 9480 11027 9482
rect 10133 9424 10138 9480
rect 10194 9424 10966 9480
rect 11022 9424 11027 9480
rect 10133 9422 11027 9424
rect 10133 9419 10199 9422
rect 10961 9419 11027 9422
rect 11145 9482 11211 9485
rect 11286 9482 11346 9694
rect 11421 9691 11487 9694
rect 15561 9618 15627 9621
rect 19600 9618 20000 9648
rect 15561 9616 20000 9618
rect 15561 9560 15566 9616
rect 15622 9560 20000 9616
rect 15561 9558 20000 9560
rect 15561 9555 15627 9558
rect 19600 9528 20000 9558
rect 11145 9480 11346 9482
rect 11145 9424 11150 9480
rect 11206 9424 11346 9480
rect 11145 9422 11346 9424
rect 11145 9419 11211 9422
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 7833 8938 7899 8941
rect 9622 8938 9628 8940
rect 7833 8936 9628 8938
rect 7833 8880 7838 8936
rect 7894 8880 9628 8936
rect 7833 8878 9628 8880
rect 7833 8875 7899 8878
rect 9622 8876 9628 8878
rect 9692 8876 9698 8940
rect 9857 8938 9923 8941
rect 10501 8938 10567 8941
rect 12893 8938 12959 8941
rect 9857 8936 12959 8938
rect 9857 8880 9862 8936
rect 9918 8880 10506 8936
rect 10562 8880 12898 8936
rect 12954 8880 12959 8936
rect 9857 8878 12959 8880
rect 9857 8875 9923 8878
rect 10501 8875 10567 8878
rect 12893 8875 12959 8878
rect 19057 8938 19123 8941
rect 19600 8938 20000 8968
rect 19057 8936 20000 8938
rect 19057 8880 19062 8936
rect 19118 8880 20000 8936
rect 19057 8878 20000 8880
rect 19057 8875 19123 8878
rect 19600 8848 20000 8878
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 11145 8530 11211 8533
rect 12525 8530 12591 8533
rect 11145 8528 12591 8530
rect 11145 8472 11150 8528
rect 11206 8472 12530 8528
rect 12586 8472 12591 8528
rect 11145 8470 12591 8472
rect 11145 8467 11211 8470
rect 12525 8467 12591 8470
rect 11697 8258 11763 8261
rect 12157 8258 12223 8261
rect 11697 8256 12223 8258
rect 11697 8200 11702 8256
rect 11758 8200 12162 8256
rect 12218 8200 12223 8256
rect 11697 8198 12223 8200
rect 11697 8195 11763 8198
rect 12157 8195 12223 8198
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19600 8168 20000 8288
rect 19253 8127 19569 8128
rect 11513 8122 11579 8125
rect 12985 8122 13051 8125
rect 11513 8120 13051 8122
rect 11513 8064 11518 8120
rect 11574 8064 12990 8120
rect 13046 8064 13051 8120
rect 11513 8062 13051 8064
rect 11513 8059 11579 8062
rect 12985 8059 13051 8062
rect 12433 7986 12499 7989
rect 13721 7986 13787 7989
rect 12433 7984 13787 7986
rect 12433 7928 12438 7984
rect 12494 7928 13726 7984
rect 13782 7928 13787 7984
rect 12433 7926 13787 7928
rect 12433 7923 12499 7926
rect 13721 7923 13787 7926
rect 19750 7853 19810 8168
rect 12433 7850 12499 7853
rect 12893 7850 12959 7853
rect 12433 7848 12959 7850
rect 12433 7792 12438 7848
rect 12494 7792 12898 7848
rect 12954 7792 12959 7848
rect 12433 7790 12959 7792
rect 12433 7787 12499 7790
rect 12893 7787 12959 7790
rect 19701 7848 19810 7853
rect 19701 7792 19706 7848
rect 19762 7792 19810 7848
rect 19701 7790 19810 7792
rect 19701 7787 19767 7790
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 19057 7578 19123 7581
rect 19600 7578 20000 7608
rect 19057 7576 20000 7578
rect 19057 7520 19062 7576
rect 19118 7520 20000 7576
rect 19057 7518 20000 7520
rect 19057 7515 19123 7518
rect 19600 7488 20000 7518
rect 11697 7442 11763 7445
rect 13905 7442 13971 7445
rect 11697 7440 13971 7442
rect 11697 7384 11702 7440
rect 11758 7384 13910 7440
rect 13966 7384 13971 7440
rect 11697 7382 13971 7384
rect 11697 7379 11763 7382
rect 13905 7379 13971 7382
rect 13721 7306 13787 7309
rect 16665 7306 16731 7309
rect 13721 7304 16731 7306
rect 13721 7248 13726 7304
rect 13782 7248 16670 7304
rect 16726 7248 16731 7304
rect 13721 7246 16731 7248
rect 13721 7243 13787 7246
rect 16665 7243 16731 7246
rect 13629 7170 13695 7173
rect 13997 7170 14063 7173
rect 13629 7168 14063 7170
rect 13629 7112 13634 7168
rect 13690 7112 14002 7168
rect 14058 7112 14063 7168
rect 13629 7110 14063 7112
rect 13629 7107 13695 7110
rect 13997 7107 14063 7110
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 15193 6898 15259 6901
rect 16849 6898 16915 6901
rect 15193 6896 16915 6898
rect 15193 6840 15198 6896
rect 15254 6840 16854 6896
rect 16910 6840 16915 6896
rect 15193 6838 16915 6840
rect 15193 6835 15259 6838
rect 16849 6835 16915 6838
rect 19425 6898 19491 6901
rect 19600 6898 20000 6928
rect 19425 6896 20000 6898
rect 19425 6840 19430 6896
rect 19486 6840 20000 6896
rect 19425 6838 20000 6840
rect 19425 6835 19491 6838
rect 19600 6808 20000 6838
rect 13721 6762 13787 6765
rect 14917 6762 14983 6765
rect 17401 6762 17467 6765
rect 13721 6760 17467 6762
rect 13721 6704 13726 6760
rect 13782 6704 14922 6760
rect 14978 6704 17406 6760
rect 17462 6704 17467 6760
rect 13721 6702 17467 6704
rect 13721 6699 13787 6702
rect 14917 6699 14983 6702
rect 17401 6699 17467 6702
rect 12801 6626 12867 6629
rect 14273 6626 14339 6629
rect 12801 6624 14339 6626
rect 12801 6568 12806 6624
rect 12862 6568 14278 6624
rect 14334 6568 14339 6624
rect 12801 6566 14339 6568
rect 12801 6563 12867 6566
rect 14273 6563 14339 6566
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 4337 6354 4403 6357
rect 5165 6354 5231 6357
rect 4337 6352 5231 6354
rect 4337 6296 4342 6352
rect 4398 6296 5170 6352
rect 5226 6296 5231 6352
rect 4337 6294 5231 6296
rect 4337 6291 4403 6294
rect 5165 6291 5231 6294
rect 13169 6354 13235 6357
rect 15653 6354 15719 6357
rect 13169 6352 15719 6354
rect 13169 6296 13174 6352
rect 13230 6296 15658 6352
rect 15714 6296 15719 6352
rect 13169 6294 15719 6296
rect 13169 6291 13235 6294
rect 15653 6291 15719 6294
rect 4613 6218 4679 6221
rect 5441 6218 5507 6221
rect 4613 6216 5507 6218
rect 4613 6160 4618 6216
rect 4674 6160 5446 6216
rect 5502 6160 5507 6216
rect 4613 6158 5507 6160
rect 4613 6155 4679 6158
rect 5441 6155 5507 6158
rect 13353 6218 13419 6221
rect 14089 6218 14155 6221
rect 13353 6216 14155 6218
rect 13353 6160 13358 6216
rect 13414 6160 14094 6216
rect 14150 6160 14155 6216
rect 13353 6158 14155 6160
rect 13353 6155 13419 6158
rect 14089 6155 14155 6158
rect 18689 6218 18755 6221
rect 19600 6218 20000 6248
rect 18689 6216 20000 6218
rect 18689 6160 18694 6216
rect 18750 6160 20000 6216
rect 18689 6158 20000 6160
rect 18689 6155 18755 6158
rect 19600 6128 20000 6158
rect 12985 6082 13051 6085
rect 13629 6082 13695 6085
rect 12985 6080 13695 6082
rect 12985 6024 12990 6080
rect 13046 6024 13634 6080
rect 13690 6024 13695 6080
rect 12985 6022 13695 6024
rect 12985 6019 13051 6022
rect 13629 6019 13695 6022
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 11421 5946 11487 5949
rect 12566 5946 12572 5948
rect 11421 5944 12572 5946
rect 11421 5888 11426 5944
rect 11482 5888 12572 5944
rect 11421 5886 12572 5888
rect 11421 5883 11487 5886
rect 12566 5884 12572 5886
rect 12636 5884 12642 5948
rect 16297 5810 16363 5813
rect 15150 5808 16363 5810
rect 15150 5752 16302 5808
rect 16358 5752 16363 5808
rect 15150 5750 16363 5752
rect 15150 5677 15210 5750
rect 16297 5747 16363 5750
rect 12341 5674 12407 5677
rect 15101 5674 15210 5677
rect 12341 5672 15210 5674
rect 12341 5616 12346 5672
rect 12402 5616 15106 5672
rect 15162 5616 15210 5672
rect 12341 5614 15210 5616
rect 15285 5674 15351 5677
rect 18781 5674 18847 5677
rect 15285 5672 18847 5674
rect 15285 5616 15290 5672
rect 15346 5616 18786 5672
rect 18842 5616 18847 5672
rect 15285 5614 18847 5616
rect 12341 5611 12407 5614
rect 15101 5611 15167 5614
rect 15285 5611 15351 5614
rect 18781 5611 18847 5614
rect 15377 5538 15443 5541
rect 16389 5538 16455 5541
rect 15377 5536 16455 5538
rect 15377 5480 15382 5536
rect 15438 5480 16394 5536
rect 16450 5480 16455 5536
rect 15377 5478 16455 5480
rect 15377 5475 15443 5478
rect 16389 5475 16455 5478
rect 18597 5538 18663 5541
rect 19600 5538 20000 5568
rect 18597 5536 20000 5538
rect 18597 5480 18602 5536
rect 18658 5480 20000 5536
rect 18597 5478 20000 5480
rect 18597 5475 18663 5478
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 19600 5448 20000 5478
rect 16896 5407 17212 5408
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 0 4178 400 4208
rect 473 4178 539 4181
rect 0 4176 539 4178
rect 0 4120 478 4176
rect 534 4120 539 4176
rect 0 4118 539 4120
rect 0 4088 400 4118
rect 473 4115 539 4118
rect 8477 4178 8543 4181
rect 15469 4178 15535 4181
rect 8477 4176 15535 4178
rect 8477 4120 8482 4176
rect 8538 4120 15474 4176
rect 15530 4120 15535 4176
rect 8477 4118 15535 4120
rect 8477 4115 8543 4118
rect 15469 4115 15535 4118
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19600 2728 20000 2848
rect 19253 2687 19569 2688
rect 19609 2410 19675 2413
rect 19750 2410 19810 2728
rect 19609 2408 19810 2410
rect 19609 2352 19614 2408
rect 19670 2352 19810 2408
rect 19609 2350 19810 2352
rect 19609 2347 19675 2350
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 19057 2138 19123 2141
rect 19600 2138 20000 2168
rect 19057 2136 20000 2138
rect 19057 2080 19062 2136
rect 19118 2080 20000 2136
rect 19057 2078 20000 2080
rect 19057 2075 19123 2078
rect 19600 2048 20000 2078
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 0 1458 400 1488
rect 841 1458 907 1461
rect 0 1456 907 1458
rect 0 1400 846 1456
rect 902 1400 907 1456
rect 0 1398 907 1400
rect 0 1368 400 1398
rect 841 1395 907 1398
rect 18873 1458 18939 1461
rect 19600 1458 20000 1488
rect 18873 1456 20000 1458
rect 18873 1400 18878 1456
rect 18934 1400 20000 1456
rect 18873 1398 20000 1400
rect 18873 1395 18939 1398
rect 19600 1368 20000 1398
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 9260 15268 9324 15332
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 9628 12820 9692 12884
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 12572 11052 12636 11116
rect 9260 10916 9324 10980
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 9628 8876 9692 8940
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 12572 5884 12636 5948
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 9259 15332 9325 15333
rect 9259 15268 9260 15332
rect 9324 15268 9325 15332
rect 9259 15267 9325 15268
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 9262 10981 9322 15267
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 9627 12884 9693 12885
rect 9627 12820 9628 12884
rect 9692 12820 9693 12884
rect 9627 12819 9693 12820
rect 9259 10980 9325 10981
rect 9259 10916 9260 10980
rect 9324 10916 9325 10980
rect 9259 10915 9325 10916
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 9630 8941 9690 12819
rect 9821 12544 10141 13568
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 9821 11456 10141 12480
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9627 8940 9693 8941
rect 9627 8876 9628 8940
rect 9692 8876 9693 8940
rect 9627 8875 9693 8876
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 12571 11116 12637 11117
rect 12571 11052 12572 11116
rect 12636 11052 12637 11116
rect 12571 11051 12637 11052
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 12179 5472 12499 6496
rect 12574 5949 12634 11051
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 12571 5948 12637 5949
rect 12571 5884 12572 5948
rect 12636 5884 12637 5948
rect 12571 5883 12637 5884
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 12179 496 12499 1056
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__nor2_2  _241_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 8832 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _242_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8464 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _243_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 8740 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _244_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8740 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _245_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _246_
timestamp 1701704242
transform -1 0 11776 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _247_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9568 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _248_
timestamp 1701704242
transform -1 0 12512 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1701704242
transform -1 0 8280 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _250_
timestamp 1701704242
transform -1 0 12328 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1701704242
transform -1 0 8188 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _252_
timestamp 1701704242
transform -1 0 8740 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _253_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _254_
timestamp 1701704242
transform -1 0 10396 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _255_
timestamp 1701704242
transform -1 0 12512 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _256_
timestamp 1701704242
transform -1 0 10580 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _257_
timestamp 1701704242
transform -1 0 11316 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _258_
timestamp 1701704242
transform -1 0 10856 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _259_
timestamp 1701704242
transform 1 0 9016 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__or3b_2  _260_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12420 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _261_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16008 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _262_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16560 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _263_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1701704242
transform -1 0 13800 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _265_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _266_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14260 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _267_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13524 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _268_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _269_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16008 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _270_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17388 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _271_
timestamp 1701704242
transform -1 0 16560 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _272_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16468 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _273_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _274_
timestamp 1701704242
transform -1 0 16376 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _275_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12604 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _276_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15272 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _277_
timestamp 1701704242
transform -1 0 15824 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _278_
timestamp 1701704242
transform -1 0 16928 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _279_
timestamp 1701704242
transform -1 0 17480 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _280_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15456 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _281_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10396 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _282_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14628 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _283_
timestamp 1701704242
transform -1 0 13984 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _284_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12512 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _285_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _286_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13892 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _287_
timestamp 1701704242
transform -1 0 14444 0 -1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_2  _288_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14352 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _289_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12512 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _290_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7820 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _291_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _292_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13248 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _293_
timestamp 1701704242
transform -1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _294_
timestamp 1701704242
transform -1 0 13800 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _295_
timestamp 1701704242
transform -1 0 14444 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _296_
timestamp 1701704242
transform -1 0 10396 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _297_
timestamp 1701704242
transform 1 0 9476 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _298_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_2  _299_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15916 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_2  _300_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15640 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_2  _301_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18216 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_4  _302_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12512 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_4  _303_
timestamp 1701704242
transform -1 0 17480 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _304_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15916 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _305_
timestamp 1701704242
transform -1 0 11960 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _306_
timestamp 1701704242
transform 1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _307_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _308_
timestamp 1701704242
transform 1 0 12696 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _309_
timestamp 1701704242
transform 1 0 11868 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _310_
timestamp 1701704242
transform 1 0 12236 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _311_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11408 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _312_
timestamp 1701704242
transform 1 0 11684 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp 1701704242
transform 1 0 8464 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _314_
timestamp 1701704242
transform 1 0 10212 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _315_
timestamp 1701704242
transform 1 0 12420 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_4  _316_
timestamp 1701704242
transform -1 0 15640 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ai_4  _317_
timestamp 1701704242
transform -1 0 17296 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _318_
timestamp 1701704242
transform 1 0 11132 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _319_
timestamp 1701704242
transform 1 0 11684 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _320_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _321_
timestamp 1701704242
transform -1 0 16008 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _322_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12236 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _323_
timestamp 1701704242
transform -1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _324_
timestamp 1701704242
transform -1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _325_
timestamp 1701704242
transform -1 0 12236 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _326_
timestamp 1701704242
transform 1 0 10580 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _327_
timestamp 1701704242
transform 1 0 10212 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _328_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11316 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _329_
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _330_
timestamp 1701704242
transform 1 0 11132 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _331_
timestamp 1701704242
transform 1 0 12604 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _332_
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _333_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12052 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _334_
timestamp 1701704242
transform 1 0 12052 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_4  _335_
timestamp 1701704242
transform -1 0 13432 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_2  _336_
timestamp 1701704242
transform -1 0 18216 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _337_
timestamp 1701704242
transform 1 0 10120 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _338_
timestamp 1701704242
transform -1 0 10764 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _339_
timestamp 1701704242
transform -1 0 11592 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1701704242
transform 1 0 7176 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _341_
timestamp 1701704242
transform -1 0 9568 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _342_
timestamp 1701704242
transform 1 0 7820 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _343_
timestamp 1701704242
transform 1 0 8556 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _344_
timestamp 1701704242
transform 1 0 9568 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _345_
timestamp 1701704242
transform 1 0 15640 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _346_
timestamp 1701704242
transform 1 0 13984 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _347_
timestamp 1701704242
transform -1 0 12052 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _348_
timestamp 1701704242
transform -1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _349_
timestamp 1701704242
transform 1 0 5152 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _350_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14168 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__a31o_1  _351_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13156 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _352_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _353_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16928 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _354_
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _355_
timestamp 1701704242
transform -1 0 19044 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_4  _356_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13156 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _357_
timestamp 1701704242
transform 1 0 18216 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _358_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12696 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _359_
timestamp 1701704242
transform 1 0 8096 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _360_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15456 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_8  _361_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15272 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_1  _362_
timestamp 1701704242
transform 1 0 13248 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 1701704242
transform 1 0 11408 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _364_
timestamp 1701704242
transform 1 0 15916 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _365_
timestamp 1701704242
transform -1 0 19136 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _366_
timestamp 1701704242
transform -1 0 18216 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _367_
timestamp 1701704242
transform -1 0 19136 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _368_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _369_
timestamp 1701704242
transform 1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _370_
timestamp 1701704242
transform -1 0 17480 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _371_
timestamp 1701704242
transform -1 0 19136 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _372_
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _373_
timestamp 1701704242
transform 1 0 17388 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _374_
timestamp 1701704242
transform -1 0 19136 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _375_
timestamp 1701704242
transform -1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376__1
timestamp 1701704242
transform 1 0 2852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377__2
timestamp 1701704242
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _378_
timestamp 1701704242
transform -1 0 11408 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _379_
timestamp 1701704242
transform -1 0 9752 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _380_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10304 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _381_
timestamp 1701704242
transform 1 0 9844 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _382_
timestamp 1701704242
transform -1 0 11408 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _383_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 11776 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _384_
timestamp 1701704242
transform -1 0 16652 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _385__3
timestamp 1701704242
transform -1 0 8280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386__4
timestamp 1701704242
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1701704242
transform 1 0 9936 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1701704242
transform -1 0 9752 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _389_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10028 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _390_
timestamp 1701704242
transform 1 0 10120 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _391_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10028 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _392_
timestamp 1701704242
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _393_
timestamp 1701704242
transform 1 0 1472 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _394_
timestamp 1701704242
transform -1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _395_
timestamp 1701704242
transform -1 0 3128 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp 1701704242
transform 1 0 2392 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _397_
timestamp 1701704242
transform -1 0 3588 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _398_
timestamp 1701704242
transform -1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _399_
timestamp 1701704242
transform 1 0 1472 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _400_
timestamp 1701704242
transform 1 0 1288 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _401_
timestamp 1701704242
transform -1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _402_
timestamp 1701704242
transform -1 0 2760 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _403_
timestamp 1701704242
transform -1 0 2024 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _404_
timestamp 1701704242
transform 1 0 2668 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _405_
timestamp 1701704242
transform 1 0 2760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _406_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _407_
timestamp 1701704242
transform -1 0 3036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _408_
timestamp 1701704242
transform 1 0 2760 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _409_
timestamp 1701704242
transform 1 0 3404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _410_
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _411_
timestamp 1701704242
transform -1 0 3680 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _412_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _413_
timestamp 1701704242
transform -1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _414_
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _415_
timestamp 1701704242
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _416_
timestamp 1701704242
transform 1 0 4232 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _417_
timestamp 1701704242
transform -1 0 4876 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1701704242
transform -1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _419_
timestamp 1701704242
transform 1 0 3864 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _420_
timestamp 1701704242
transform -1 0 4048 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _421_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _422_
timestamp 1701704242
transform 1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _423_
timestamp 1701704242
transform 1 0 4416 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _424_
timestamp 1701704242
transform -1 0 7728 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _425_
timestamp 1701704242
transform -1 0 6992 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _426_
timestamp 1701704242
transform -1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _427_
timestamp 1701704242
transform -1 0 7544 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _428_
timestamp 1701704242
transform -1 0 6624 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _429_
timestamp 1701704242
transform -1 0 7360 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _430_
timestamp 1701704242
transform -1 0 7268 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _431_
timestamp 1701704242
transform -1 0 6992 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _432_
timestamp 1701704242
transform -1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _433_
timestamp 1701704242
transform 1 0 6348 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1701704242
transform -1 0 6624 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _435_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 6348 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _436_
timestamp 1701704242
transform 1 0 5060 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _437_
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _438_
timestamp 1701704242
transform -1 0 6256 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _439_
timestamp 1701704242
transform 1 0 4600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _440_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 4600 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _441_
timestamp 1701704242
transform -1 0 3864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _442_
timestamp 1701704242
transform 1 0 3772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _443_
timestamp 1701704242
transform 1 0 3864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _444_
timestamp 1701704242
transform -1 0 3864 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _446_
timestamp 1701704242
transform 1 0 4048 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _447_
timestamp 1701704242
transform 1 0 5152 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _448_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1701704242
transform -1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_1  _450_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4508 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _451_
timestamp 1701704242
transform 1 0 4876 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1701704242
transform -1 0 9384 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 1701704242
transform 1 0 9936 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1701704242
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _455_
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1701704242
transform 1 0 6716 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 1701704242
transform -1 0 5704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1701704242
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1701704242
transform -1 0 5612 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp 1701704242
transform 1 0 4876 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _461_
timestamp 1701704242
transform 1 0 4968 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1701704242
transform 1 0 7176 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _463_
timestamp 1701704242
transform 1 0 6992 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1701704242
transform 1 0 9384 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _465_
timestamp 1701704242
transform 1 0 9568 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1701704242
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp 1701704242
transform 1 0 6256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1701704242
transform 1 0 6164 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1701704242
transform 1 0 4968 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _470_
timestamp 1701704242
transform -1 0 8280 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp 1701704242
transform 1 0 11684 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _472_
timestamp 1701704242
transform -1 0 11592 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1701704242
transform -1 0 12512 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _474_
timestamp 1701704242
transform 1 0 12512 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1701704242
transform 1 0 8556 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp 1701704242
transform -1 0 9016 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1701704242
transform -1 0 9844 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp 1701704242
transform -1 0 10120 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 1701704242
transform 1 0 11408 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp 1701704242
transform -1 0 11224 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1701704242
transform 1 0 9936 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1701704242
transform -1 0 9844 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _484_
timestamp 1701704242
transform -1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _486_
timestamp 1701704242
transform 1 0 6440 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _487_
timestamp 1701704242
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _488_
timestamp 1701704242
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _489_
timestamp 1701704242
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _490_
timestamp 1701704242
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _492_
timestamp 1701704242
transform 1 0 6716 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _493_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1701704242
transform 1 0 1380 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _495_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _496_
timestamp 1701704242
transform 1 0 11776 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _497_
timestamp 1701704242
transform 1 0 13064 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1701704242
transform 1 0 7728 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1701704242
transform 1 0 9384 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _500_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8740 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1701704242
transform 1 0 9752 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _502_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _505_
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1701704242
transform 1 0 3128 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1701704242
transform 1 0 2852 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _508_
timestamp 1701704242
transform 1 0 2300 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _509_
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _510_
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _511_
timestamp 1701704242
transform 1 0 3588 0 -1 17952
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _512_
timestamp 1701704242
transform 1 0 6348 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _513_
timestamp 1701704242
transform 1 0 7176 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1701704242
transform 1 0 6072 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _515_
timestamp 1701704242
transform 1 0 4968 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _517_
timestamp 1701704242
transform 1 0 2208 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1701704242
transform 1 0 3404 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1701704242
transform 1 0 3864 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1701704242
transform -1 0 9936 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _521_
timestamp 1701704242
transform 1 0 7636 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _523_
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1701704242
transform 1 0 4232 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1701704242
transform 1 0 6532 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1701704242
transform 1 0 9108 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp 1701704242
transform 1 0 5796 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp 1701704242
transform 1 0 11592 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp 1701704242
transform 1 0 11684 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _531_
timestamp 1701704242
transform 1 0 9016 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 1701704242
transform -1 0 10856 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _533_
timestamp 1701704242
transform 1 0 11224 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 1701704242
transform 1 0 9844 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _535_
timestamp 1701704242
transform 1 0 7912 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 1701704242
transform 1 0 5980 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _537_
timestamp 1701704242
transform 1 0 5980 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _538_
timestamp 1701704242
transform 1 0 5980 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _539_
timestamp 1701704242
transform 1 0 6256 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7176 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1701704242
transform 1 0 4876 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1701704242
transform 1 0 7912 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1701704242
transform -1 0 6256 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1701704242
transform 1 0 7728 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  fanout1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18216 0 1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout2
timestamp 1701704242
transform -1 0 14076 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout3
timestamp 1701704242
transform 1 0 18124 0 -1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout4
timestamp 1701704242
transform -1 0 18400 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout14 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 17756 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout15
timestamp 1701704242
transform -1 0 12420 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1701704242
transform -1 0 5888 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1701704242
transform 1 0 6532 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1701704242
transform -1 0 4600 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1701704242
transform -1 0 4968 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_40
timestamp 1701704242
transform 1 0 4232 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_52 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5336 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_116 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11224 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_159
timestamp 1701704242
transform 1 0 15180 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1701704242
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_190 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18032 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_51
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_124
timestamp 1701704242
transform 1 0 11960 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_190
timestamp 1701704242
transform 1 0 18032 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_198
timestamp 1701704242
transform 1 0 18768 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 1701704242
transform 1 0 1104 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18
timestamp 1701704242
transform 1 0 2208 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1701704242
transform 1 0 2944 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_147
timestamp 1701704242
transform 1 0 14076 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_172
timestamp 1701704242
transform 1 0 16376 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_176
timestamp 1701704242
transform 1 0 16744 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_200
timestamp 1701704242
transform 1 0 18952 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_187
timestamp 1701704242
transform 1 0 17756 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_71
timestamp 1701704242
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_79
timestamp 1701704242
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_36
timestamp 1701704242
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1701704242
transform 1 0 4968 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1701704242
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_70
timestamp 1701704242
transform 1 0 6992 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_181
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_186
timestamp 1701704242
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_190
timestamp 1701704242
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_45
timestamp 1701704242
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_57
timestamp 1701704242
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_61
timestamp 1701704242
transform 1 0 6164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1701704242
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_100
timestamp 1701704242
transform 1 0 9752 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_144
timestamp 1701704242
transform 1 0 13800 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1701704242
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 1701704242
transform 1 0 1104 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 1701704242
transform 1 0 2208 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_30
timestamp 1701704242
transform 1 0 3312 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_79
timestamp 1701704242
transform 1 0 7820 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_145
timestamp 1701704242
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1701704242
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_175
timestamp 1701704242
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_51
timestamp 1701704242
transform 1 0 5244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_58
timestamp 1701704242
transform 1 0 5888 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_67
timestamp 1701704242
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_109
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_147
timestamp 1701704242
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1701704242
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_74
timestamp 1701704242
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_100
timestamp 1701704242
transform 1 0 9752 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_136
timestamp 1701704242
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_37
timestamp 1701704242
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_57
timestamp 1701704242
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_63
timestamp 1701704242
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_67
timestamp 1701704242
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1701704242
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_88
timestamp 1701704242
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_98
timestamp 1701704242
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_125
timestamp 1701704242
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1701704242
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_9
timestamp 1701704242
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_16
timestamp 1701704242
transform 1 0 2024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_30
timestamp 1701704242
transform 1 0 3312 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_79
timestamp 1701704242
transform 1 0 7820 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_100
timestamp 1701704242
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_107
timestamp 1701704242
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1701704242
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_139
timestamp 1701704242
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_149
timestamp 1701704242
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_182
timestamp 1701704242
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_24
timestamp 1701704242
transform 1 0 2760 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1701704242
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_92
timestamp 1701704242
transform 1 0 9016 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_98
timestamp 1701704242
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_103
timestamp 1701704242
transform 1 0 10028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_114
timestamp 1701704242
transform 1 0 11040 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_11
timestamp 1701704242
transform 1 0 1564 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_16
timestamp 1701704242
transform 1 0 2024 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_28
timestamp 1701704242
transform 1 0 3128 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_40
timestamp 1701704242
transform 1 0 4232 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_52
timestamp 1701704242
transform 1 0 5336 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_77
timestamp 1701704242
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1701704242
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1701704242
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_154
timestamp 1701704242
transform 1 0 14720 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_17
timestamp 1701704242
transform 1 0 2116 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1701704242
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_49
timestamp 1701704242
transform 1 0 5060 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_55
timestamp 1701704242
transform 1 0 5612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_73
timestamp 1701704242
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_98
timestamp 1701704242
transform 1 0 9568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_110
timestamp 1701704242
transform 1 0 10672 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_136
timestamp 1701704242
transform 1 0 13064 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_28
timestamp 1701704242
transform 1 0 3128 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_36
timestamp 1701704242
transform 1 0 3864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_48
timestamp 1701704242
transform 1 0 4968 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_77
timestamp 1701704242
transform 1 0 7636 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_89
timestamp 1701704242
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_97
timestamp 1701704242
transform 1 0 9476 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_107
timestamp 1701704242
transform 1 0 10396 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1701704242
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_123
timestamp 1701704242
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_135
timestamp 1701704242
transform 1 0 12972 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1701704242
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_19
timestamp 1701704242
transform 1 0 2300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1701704242
transform 1 0 2852 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_33
timestamp 1701704242
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_45
timestamp 1701704242
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_57
timestamp 1701704242
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1701704242
transform 1 0 7820 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1701704242
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_94
timestamp 1701704242
transform 1 0 9200 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_120
timestamp 1701704242
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_134
timestamp 1701704242
transform 1 0 12880 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_141
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_147
timestamp 1701704242
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_166
timestamp 1701704242
transform 1 0 15824 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1701704242
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_23
timestamp 1701704242
transform 1 0 2668 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_35
timestamp 1701704242
transform 1 0 3772 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1701704242
transform 1 0 4876 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_63
timestamp 1701704242
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_67
timestamp 1701704242
transform 1 0 6716 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_71
timestamp 1701704242
transform 1 0 7084 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_103
timestamp 1701704242
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1701704242
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_118
timestamp 1701704242
transform 1 0 11408 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_124
timestamp 1701704242
transform 1 0 11960 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_144
timestamp 1701704242
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_154
timestamp 1701704242
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1701704242
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_174
timestamp 1701704242
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_201
timestamp 1701704242
transform 1 0 19044 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1701704242
transform 1 0 1196 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_14
timestamp 1701704242
transform 1 0 1840 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1701704242
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_33
timestamp 1701704242
transform 1 0 3588 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_39
timestamp 1701704242
transform 1 0 4140 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_60
timestamp 1701704242
transform 1 0 6072 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_72
timestamp 1701704242
transform 1 0 7176 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_107
timestamp 1701704242
transform 1 0 10396 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_117
timestamp 1701704242
transform 1 0 11316 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_129
timestamp 1701704242
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1701704242
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_151
timestamp 1701704242
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_200
timestamp 1701704242
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_24
timestamp 1701704242
transform 1 0 2760 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_45
timestamp 1701704242
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_63
timestamp 1701704242
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_73
timestamp 1701704242
transform 1 0 7268 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_79
timestamp 1701704242
transform 1 0 7820 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1701704242
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_162
timestamp 1701704242
transform 1 0 15456 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1701704242
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_14
timestamp 1701704242
transform 1 0 1840 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_22
timestamp 1701704242
transform 1 0 2576 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_37
timestamp 1701704242
transform 1 0 3956 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_51
timestamp 1701704242
transform 1 0 5244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1701704242
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_91
timestamp 1701704242
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_107
timestamp 1701704242
transform 1 0 10396 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_113
timestamp 1701704242
transform 1 0 10948 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_128
timestamp 1701704242
transform 1 0 12328 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_184
timestamp 1701704242
transform 1 0 17480 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1701704242
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 1701704242
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_17
timestamp 1701704242
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_48
timestamp 1701704242
transform 1 0 4968 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_61
timestamp 1701704242
transform 1 0 6164 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_65
timestamp 1701704242
transform 1 0 6532 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_71
timestamp 1701704242
transform 1 0 7084 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_86
timestamp 1701704242
transform 1 0 8464 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_106
timestamp 1701704242
transform 1 0 10304 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_145
timestamp 1701704242
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_149
timestamp 1701704242
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_191
timestamp 1701704242
transform 1 0 18124 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_199
timestamp 1701704242
transform 1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_37
timestamp 1701704242
transform 1 0 3956 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_70
timestamp 1701704242
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1701704242
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_116
timestamp 1701704242
transform 1 0 11224 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_123
timestamp 1701704242
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1701704242
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1701704242
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1701704242
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_11
timestamp 1701704242
transform 1 0 1564 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_16
timestamp 1701704242
transform 1 0 2024 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_28
timestamp 1701704242
transform 1 0 3128 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_62
timestamp 1701704242
transform 1 0 6256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_130
timestamp 1701704242
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_140
timestamp 1701704242
transform 1 0 13432 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_187
timestamp 1701704242
transform 1 0 17756 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_197
timestamp 1701704242
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_201
timestamp 1701704242
transform 1 0 19044 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_21
timestamp 1701704242
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 1701704242
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_34
timestamp 1701704242
transform 1 0 3680 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_62
timestamp 1701704242
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_73
timestamp 1701704242
transform 1 0 7268 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1701704242
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_93
timestamp 1701704242
transform 1 0 9108 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_117
timestamp 1701704242
transform 1 0 11316 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_130
timestamp 1701704242
transform 1 0 12512 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1701704242
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_149
timestamp 1701704242
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_47
timestamp 1701704242
transform 1 0 4876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_66
timestamp 1701704242
transform 1 0 6624 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_101
timestamp 1701704242
transform 1 0 9844 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1701704242
transform 1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_130
timestamp 1701704242
transform 1 0 12512 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_142
timestamp 1701704242
transform 1 0 13616 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_160
timestamp 1701704242
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1701704242
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1701704242
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_33
timestamp 1701704242
transform 1 0 3588 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_47
timestamp 1701704242
transform 1 0 4876 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_73
timestamp 1701704242
transform 1 0 7268 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_91
timestamp 1701704242
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_113
timestamp 1701704242
transform 1 0 10948 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1701704242
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_38
timestamp 1701704242
transform 1 0 4048 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_42
timestamp 1701704242
transform 1 0 4416 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_48
timestamp 1701704242
transform 1 0 4968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_100
timestamp 1701704242
transform 1 0 9752 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 1701704242
transform 1 0 13524 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 1701704242
transform 1 0 14628 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1701704242
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_49
timestamp 1701704242
transform 1 0 5060 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_61
timestamp 1701704242
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1701704242
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_94
timestamp 1701704242
transform 1 0 9200 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1701704242
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1701704242
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1701704242
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_31
timestamp 1701704242
transform 1 0 3404 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_35
timestamp 1701704242
transform 1 0 3772 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_47
timestamp 1701704242
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_76
timestamp 1701704242
transform 1 0 7544 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_84
timestamp 1701704242
transform 1 0 8280 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_96
timestamp 1701704242
transform 1 0 9384 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1701704242
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_193
timestamp 1701704242
transform 1 0 18308 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_197
timestamp 1701704242
transform 1 0 18676 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_52
timestamp 1701704242
transform 1 0 5336 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_58
timestamp 1701704242
transform 1 0 5888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_78
timestamp 1701704242
transform 1 0 7728 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_112
timestamp 1701704242
transform 1 0 10856 0 1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_127
timestamp 1701704242
transform 1 0 12236 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1701704242
transform 1 0 19044 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_70
timestamp 1701704242
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_104
timestamp 1701704242
transform 1 0 10120 0 -1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_136
timestamp 1701704242
transform 1 0 13064 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_148
timestamp 1701704242
transform 1 0 14168 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_160
timestamp 1701704242
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_201
timestamp 1701704242
transform 1 0 19044 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_61
timestamp 1701704242
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_91
timestamp 1701704242
transform 1 0 8924 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_112
timestamp 1701704242
transform 1 0 10856 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_124
timestamp 1701704242
transform 1 0 11960 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1701704242
transform 1 0 13064 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1701704242
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_6
timestamp 1701704242
transform 1 0 1104 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_18
timestamp 1701704242
transform 1 0 2208 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_26
timestamp 1701704242
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_40
timestamp 1701704242
transform 1 0 4232 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 1701704242
transform 1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_91
timestamp 1701704242
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_101
timestamp 1701704242
transform 1 0 9844 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1701704242
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_161
timestamp 1701704242
transform 1 0 15364 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1701704242
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_173
timestamp 1701704242
transform 1 0 16468 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_185
timestamp 1701704242
transform 1 0 17572 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_194
timestamp 1701704242
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1701704242
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1701704242
transform -1 0 11684 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1701704242
transform -1 0 7268 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1701704242
transform -1 0 6532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1701704242
transform -1 0 2944 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1701704242
transform -1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1701704242
transform -1 0 4968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1701704242
transform -1 0 6532 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1701704242
transform -1 0 3036 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1701704242
transform 1 0 15180 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1701704242
transform -1 0 8004 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1701704242
transform -1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1701704242
transform -1 0 19136 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1701704242
transform -1 0 18952 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18216 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1701704242
transform -1 0 18492 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1701704242
transform -1 0 19136 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1701704242
transform -1 0 19136 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1701704242
transform -1 0 19136 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1701704242
transform -1 0 19136 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1701704242
transform -1 0 19044 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1701704242
transform -1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1701704242
transform -1 0 19136 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  load_slew5
timestamp 1701704242
transform 1 0 18216 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap6
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  max_cap21
timestamp 1701704242
transform -1 0 12512 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[0\].cap_22 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[0\].cap
timestamp 1701704242
transform -1 0 6072 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[1\].cap_29
timestamp 1701704242
transform -1 0 8924 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[1\].cap
timestamp 1701704242
transform 1 0 6716 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[2\].cap_30
timestamp 1701704242
transform -1 0 7728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[2\].cap
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[3\].cap_31
timestamp 1701704242
transform -1 0 6072 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[3\].cap
timestamp 1701704242
transform -1 0 5704 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[4\].cap_32
timestamp 1701704242
transform -1 0 8648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[4\].cap
timestamp 1701704242
transform 1 0 6992 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[5\].cap_33
timestamp 1701704242
transform 1 0 7176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[5\].cap
timestamp 1701704242
transform -1 0 9200 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[6\].cap_34
timestamp 1701704242
transform 1 0 6348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[6\].cap
timestamp 1701704242
transform 1 0 6348 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[7\].cap
timestamp 1701704242
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[7\].cap_35
timestamp 1701704242
transform -1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[8\].cap_36
timestamp 1701704242
transform 1 0 7728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[8\].cap
timestamp 1701704242
transform -1 0 11960 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[9\].cap_37
timestamp 1701704242
transform -1 0 7820 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[9\].cap
timestamp 1701704242
transform 1 0 6164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[10\].cap_23
timestamp 1701704242
transform -1 0 7728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[10\].cap
timestamp 1701704242
transform 1 0 7268 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[11\].cap_24
timestamp 1701704242
transform 1 0 6624 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[11\].cap
timestamp 1701704242
transform -1 0 11224 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[12\].cap_25
timestamp 1701704242
transform -1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[12\].cap
timestamp 1701704242
transform 1 0 6072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[13\].cap_26
timestamp 1701704242
transform -1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[13\].cap
timestamp 1701704242
transform 1 0 6072 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[14\].cap_27
timestamp 1701704242
transform -1 0 7544 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[14\].cap
timestamp 1701704242
transform 1 0 6440 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ts.ts_core.capload\[15\].cap
timestamp 1701704242
transform -1 0 6348 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.capload\[15\].cap_28
timestamp 1701704242
transform 1 0 5888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 17480 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 16928 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform 1 0 16928 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform -1 0 17572 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform 1 0 16560 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 16928 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform -1 0 15548 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 15548 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform 1 0 14260 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform -1 0 16836 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1701704242
transform 1 0 13892 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1701704242
transform -1 0 15916 0 -1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1701704242
transform -1 0 15180 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform -1 0 16008 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform 1 0 13708 0 -1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform -1 0 12604 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1701704242
transform 1 0 9200 0 -1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1701704242
transform 1 0 14720 0 1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1701704242
transform -1 0 10856 0 1 544
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1701704242
transform 1 0 9200 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1701704242
transform -1 0 10120 0 1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1701704242
transform 1 0 11776 0 1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1701704242
transform 1 0 12604 0 -1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1701704242
transform 1 0 10120 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1701704242
transform -1 0 13432 0 1 544
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1701704242
transform 1 0 10120 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1701704242
transform 1 0 10120 0 1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1701704242
transform 1 0 11776 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1701704242
transform -1 0 15456 0 1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1701704242
transform -1 0 13432 0 1 3808
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1701704242
transform 1 0 15272 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1701704242
transform 1 0 8464 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1701704242
transform 1 0 15456 0 1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1701704242
transform 1 0 14352 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1701704242
transform -1 0 15180 0 1 544
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1701704242
transform -1 0 18584 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1701704242
transform 1 0 7544 0 -1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1701704242
transform 1 0 17480 0 -1 15776
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1701704242
transform 1 0 16836 0 1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1701704242
transform -1 0 13432 0 1 4896
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1701704242
transform 1 0 16468 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1701704242
transform 1 0 6624 0 1 544
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1701704242
transform 1 0 16928 0 -1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1701704242
transform -1 0 16284 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1701704242
transform -1 0 16928 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1701704242
transform 1 0 17388 0 -1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1701704242
transform 1 0 15916 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1701704242
transform 1 0 16376 0 -1 1632
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1701704242
transform 1 0 16468 0 -1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1701704242
transform 1 0 14260 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1701704242
transform 1 0 16284 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1701704242
transform 1 0 17480 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1701704242
transform 1 0 16376 0 1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1701704242
transform 1 0 14352 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1701704242
transform 1 0 17480 0 -1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.dac.vdac_single.einvp_batch\[0\].pupd_47
timestamp 1701704242
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  ts.ts_core.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1701704242
transform -1 0 16928 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  ts.ts_core.dac.vdac_single.einvp_batch\[0\].vref_38
timestamp 1701704242
transform 1 0 18400 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ts.ts_core.dac.vdac_single.einvp_batch\[0\].vref pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 19136 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ts.ts_core.dcdc
timestamp 1701704242
transform 1 0 13616 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ts.ts_core.inv1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 7176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  ts.ts_core.inv2
timestamp 1701704242
transform 1 0 6348 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_39
timestamp 1701704242
transform -1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_40
timestamp 1701704242
transform -1 0 4232 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_41
timestamp 1701704242
transform -1 0 16468 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_42
timestamp 1701704242
transform 1 0 18860 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_43
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_44
timestamp 1701704242
transform 1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_45
timestamp 1701704242
transform -1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_46
timestamp 1701704242
transform -1 0 15824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_48
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_49
timestamp 1701704242
transform 1 0 17756 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_50
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tempsens_51
timestamp 1701704242
transform 1 0 3956 0 -1 19040
box -38 -48 314 592
<< labels >>
flabel metal4 s 5106 496 5426 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9821 496 10141 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14536 496 14856 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19251 496 19571 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2749 496 3069 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7464 496 7784 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12179 496 12499 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16894 496 17214 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 17688 400 17808 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 400 0 FreeSans 224 90 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 4088 400 4208 0 FreeSans 480 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 19600 7488 20000 7608 0 FreeSans 480 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 19600 8848 20000 8968 0 FreeSans 480 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 19600 5448 20000 5568 0 FreeSans 480 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 19600 6128 20000 6248 0 FreeSans 480 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 19600 6808 20000 6928 0 FreeSans 480 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 19600 8168 20000 8288 0 FreeSans 480 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal2 s 7746 19600 7802 20000 0 FreeSans 224 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 19600 12248 20000 12368 0 FreeSans 480 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 19600 12928 20000 13048 0 FreeSans 480 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 19600 14968 20000 15088 0 FreeSans 480 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 19600 14288 20000 14408 0 FreeSans 480 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 19600 13608 20000 13728 0 FreeSans 480 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal2 s 662 0 718 400 0 FreeSans 224 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal2 s 1306 0 1362 400 0 FreeSans 224 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal2 s 1950 0 2006 400 0 FreeSans 224 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal2 s 2594 0 2650 400 0 FreeSans 224 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 1368 400 1488 0 FreeSans 480 0 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal3 s 19600 2048 20000 2168 0 FreeSans 480 0 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal3 s 0 18368 400 18488 0 FreeSans 480 0 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal2 s 3882 19600 3938 20000 0 FreeSans 224 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal3 s 19600 1368 20000 1488 0 FreeSans 480 0 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal3 s 19600 2728 20000 2848 0 FreeSans 480 0 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal3 s 19600 9528 20000 9648 0 FreeSans 480 0 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal3 s 19600 10208 20000 10328 0 FreeSans 480 0 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal2 s 8390 19600 8446 20000 0 FreeSans 224 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal3 s 19600 10888 20000 11008 0 FreeSans 480 0 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal3 s 19600 11568 20000 11688 0 FreeSans 480 0 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal3 s 0 10888 400 11008 0 FreeSans 480 0 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal2 s 9678 19600 9734 20000 0 FreeSans 224 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal2 s 10322 19600 10378 20000 0 FreeSans 224 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal2 s 10966 19600 11022 20000 0 FreeSans 224 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal2 s 9034 19600 9090 20000 0 FreeSans 224 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 10061 19040 10061 19040 0 VGND
rlabel metal1 9982 18496 9982 18496 0 VPWR
rlabel metal1 11316 3638 11316 3638 0 _004_
rlabel metal1 11592 4726 11592 4726 0 _005_
rlabel metal1 14168 3502 14168 3502 0 _006_
rlabel metal1 9200 5066 9200 5066 0 _007_
rlabel metal1 10120 6290 10120 6290 0 _008_
rlabel metal1 1334 6766 1334 6766 0 _009_
rlabel metal1 1334 8602 1334 8602 0 _010_
rlabel metal1 1242 10778 1242 10778 0 _011_
rlabel metal1 1472 12818 1472 12818 0 _012_
rlabel metal2 3358 12342 3358 12342 0 _013_
rlabel metal1 3220 10778 3220 10778 0 _014_
rlabel metal2 2622 14212 2622 14212 0 _015_
rlabel metal1 1288 14586 1288 14586 0 _016_
rlabel metal1 3496 15946 3496 15946 0 _017_
rlabel metal1 4186 17306 4186 17306 0 _018_
rlabel metal2 6118 17714 6118 17714 0 _019_
rlabel metal1 7360 17306 7360 17306 0 _020_
rlabel metal2 6394 16014 6394 16014 0 _021_
rlabel metal1 5244 14858 5244 14858 0 _022_
rlabel metal1 3581 8602 3581 8602 0 _023_
rlabel metal2 2530 6222 2530 6222 0 _024_
rlabel metal1 3949 5338 3949 5338 0 _025_
rlabel metal1 4324 4726 4324 4726 0 _026_
rlabel metal1 9798 3502 9798 3502 0 _027_
rlabel metal1 8142 5678 8142 5678 0 _028_
rlabel metal1 5888 7854 5888 7854 0 _029_
rlabel metal1 5842 9078 5842 9078 0 _030_
rlabel metal1 4692 10506 4692 10506 0 _031_
rlabel metal1 6992 13430 6992 13430 0 _032_
rlabel metal1 9522 14586 9522 14586 0 _033_
rlabel metal1 6164 11730 6164 11730 0 _034_
rlabel metal1 4830 12818 4830 12818 0 _035_
rlabel metal1 11730 14858 11730 14858 0 _036_
rlabel metal2 12282 15742 12282 15742 0 _037_
rlabel metal1 9154 17034 9154 17034 0 _038_
rlabel metal1 10166 17850 10166 17850 0 _039_
rlabel metal1 11362 17782 11362 17782 0 _040_
rlabel metal1 9982 15946 9982 15946 0 _041_
rlabel metal2 8234 15368 8234 15368 0 _042_
rlabel metal1 6348 9554 6348 9554 0 _043_
rlabel metal1 6394 6426 6394 6426 0 _044_
rlabel metal1 6302 4760 6302 4760 0 _045_
rlabel metal1 6670 3706 6670 3706 0 _046_
rlabel viali 9614 13364 9614 13364 0 _047_
rlabel metal1 9154 11186 9154 11186 0 _048_
rlabel metal1 8970 11050 8970 11050 0 _049_
rlabel metal1 12650 8364 12650 8364 0 _050_
rlabel metal1 9706 11628 9706 11628 0 _051_
rlabel metal1 9292 8602 9292 8602 0 _052_
rlabel metal1 8602 8602 8602 8602 0 _053_
rlabel metal1 9430 10608 9430 10608 0 _054_
rlabel metal1 8786 9146 8786 9146 0 _055_
rlabel metal1 10236 12750 10236 12750 0 _056_
rlabel metal1 10534 13362 10534 13362 0 _057_
rlabel viali 11822 7922 11822 7922 0 _058_
rlabel metal2 14536 13158 14536 13158 0 _059_
rlabel metal2 12374 6732 12374 6732 0 _060_
rlabel metal1 13754 8364 13754 8364 0 _061_
rlabel metal2 12558 5746 12558 5746 0 _062_
rlabel metal1 12788 5270 12788 5270 0 _063_
rlabel metal1 14398 8976 14398 8976 0 _064_
rlabel metal2 15134 7344 15134 7344 0 _065_
rlabel metal2 12926 13838 12926 13838 0 _066_
rlabel metal2 15042 10370 15042 10370 0 _067_
rlabel metal2 13478 12580 13478 12580 0 _068_
rlabel metal1 11194 9044 11194 9044 0 _069_
rlabel metal1 11500 7922 11500 7922 0 _070_
rlabel metal1 10994 12818 10994 12818 0 _071_
rlabel metal2 13018 13804 13018 13804 0 _072_
rlabel metal1 15042 9894 15042 9894 0 _073_
rlabel metal1 14950 11084 14950 11084 0 _074_
rlabel metal1 9154 7922 9154 7922 0 _075_
rlabel metal1 10488 10642 10488 10642 0 _076_
rlabel metal1 13616 11186 13616 11186 0 _077_
rlabel metal1 13018 11050 13018 11050 0 _078_
rlabel metal1 11316 10778 11316 10778 0 _079_
rlabel metal1 11224 10098 11224 10098 0 _080_
rlabel via1 13215 13362 13215 13362 0 _081_
rlabel metal1 12098 13464 12098 13464 0 _082_
rlabel metal1 8234 12240 8234 12240 0 _083_
rlabel metal1 12650 12070 12650 12070 0 _084_
rlabel metal1 8326 12410 8326 12410 0 _085_
rlabel metal2 11086 10557 11086 10557 0 _086_
rlabel metal1 12742 10098 12742 10098 0 _087_
rlabel metal1 13202 12648 13202 12648 0 _088_
rlabel metal2 13294 9350 13294 9350 0 _089_
rlabel metal1 12995 10710 12995 10710 0 _090_
rlabel metal1 9936 9146 9936 9146 0 _091_
rlabel metal1 10396 9690 10396 9690 0 _092_
rlabel metal1 11546 9894 11546 9894 0 _093_
rlabel metal1 15870 8942 15870 8942 0 _094_
rlabel metal2 15410 10166 15410 10166 0 _095_
rlabel metal1 12282 7956 12282 7956 0 _096_
rlabel via1 15138 9486 15138 9486 0 _097_
rlabel metal1 13984 5746 13984 5746 0 _098_
rlabel metal2 16146 9384 16146 9384 0 _099_
rlabel metal1 14950 8942 14950 8942 0 _100_
rlabel metal1 12696 12954 12696 12954 0 _101_
rlabel metal2 12558 13056 12558 13056 0 _102_
rlabel metal2 12558 11084 12558 11084 0 _103_
rlabel metal2 11822 9248 11822 9248 0 _104_
rlabel metal1 12466 9656 12466 9656 0 _105_
rlabel metal1 9660 8058 9660 8058 0 _106_
rlabel metal1 12466 9520 12466 9520 0 _107_
rlabel metal1 14950 9044 14950 9044 0 _108_
rlabel metal2 11638 8194 11638 8194 0 _109_
rlabel metal1 12650 7242 12650 7242 0 _110_
rlabel metal1 15042 7310 15042 7310 0 _111_
rlabel metal1 13340 6834 13340 6834 0 _112_
rlabel metal1 12834 7820 12834 7820 0 _113_
rlabel metal1 13524 6630 13524 6630 0 _114_
rlabel metal1 13570 6732 13570 6732 0 _115_
rlabel metal1 11730 12410 11730 12410 0 _116_
rlabel metal1 11316 12818 11316 12818 0 _117_
rlabel metal1 11224 12750 11224 12750 0 _118_
rlabel metal1 11960 12614 11960 12614 0 _119_
rlabel metal1 11362 9520 11362 9520 0 _120_
rlabel metal1 11914 13158 11914 13158 0 _121_
rlabel metal1 12834 7922 12834 7922 0 _122_
rlabel metal1 9660 7514 9660 7514 0 _123_
rlabel metal1 12052 8330 12052 8330 0 _124_
rlabel viali 13202 7308 13202 7308 0 _125_
rlabel metal3 10672 9724 10672 9724 0 _126_
rlabel metal1 10994 9520 10994 9520 0 _127_
rlabel metal1 11270 9690 11270 9690 0 _128_
rlabel metal1 9292 10098 9292 10098 0 _129_
rlabel metal1 9568 9894 9568 9894 0 _130_
rlabel metal2 8602 12585 8602 12585 0 _131_
rlabel metal1 9384 12614 9384 12614 0 _132_
rlabel metal1 13570 9554 13570 9554 0 _133_
rlabel metal2 14490 9316 14490 9316 0 _134_
rlabel metal2 14674 9690 14674 9690 0 _135_
rlabel metal1 6394 6222 6394 6222 0 _136_
rlabel metal1 5934 14348 5934 14348 0 _137_
rlabel metal1 2024 14450 2024 14450 0 _138_
rlabel metal1 8234 4692 8234 4692 0 _139_
rlabel metal1 14582 8330 14582 8330 0 _140_
rlabel metal1 18860 6222 18860 6222 0 _141_
rlabel metal2 18906 4093 18906 4093 0 _142_
rlabel metal1 15134 7378 15134 7378 0 _143_
rlabel metal2 8326 4454 8326 4454 0 _144_
rlabel metal2 8510 4301 8510 4301 0 _145_
rlabel metal1 13616 5610 13616 5610 0 _146_
rlabel metal2 12742 5372 12742 5372 0 _147_
rlabel metal1 18538 7310 18538 7310 0 _148_
rlabel metal1 13202 8500 13202 8500 0 _149_
rlabel metal1 17664 4794 17664 4794 0 _150_
rlabel viali 13570 7311 13570 7311 0 _151_
rlabel metal2 18722 10132 18722 10132 0 _152_
rlabel metal2 9614 4930 9614 4930 0 _153_
rlabel metal2 7866 13396 7866 13396 0 _154_
rlabel metal2 10810 4318 10810 4318 0 _155_
rlabel metal1 11178 4590 11178 4590 0 _156_
rlabel metal1 9844 5746 9844 5746 0 _157_
rlabel metal1 9890 6698 9890 6698 0 _158_
rlabel metal1 9982 7378 9982 7378 0 _159_
rlabel metal2 1702 7276 1702 7276 0 _160_
rlabel metal1 1840 8534 1840 8534 0 _161_
rlabel metal2 3174 9860 3174 9860 0 _162_
rlabel metal1 3128 9418 3128 9418 0 _163_
rlabel metal2 1702 9486 1702 9486 0 _164_
rlabel metal2 1518 11186 1518 11186 0 _165_
rlabel metal1 1978 12138 1978 12138 0 _166_
rlabel metal1 2254 12070 2254 12070 0 _167_
rlabel metal2 3082 12517 3082 12517 0 _168_
rlabel metal1 2990 12206 2990 12206 0 _169_
rlabel metal2 3358 11254 3358 11254 0 _170_
rlabel metal1 3450 10098 3450 10098 0 _171_
rlabel metal1 3404 14926 3404 14926 0 _172_
rlabel metal1 2208 14450 2208 14450 0 _173_
rlabel metal1 2806 13872 2806 13872 0 _174_
rlabel metal1 1656 14450 1656 14450 0 _175_
rlabel metal1 4876 14586 4876 14586 0 _176_
rlabel metal1 4508 15538 4508 15538 0 _177_
rlabel metal1 4048 15334 4048 15334 0 _178_
rlabel metal2 3910 15368 3910 15368 0 _179_
rlabel metal1 3680 15402 3680 15402 0 _180_
rlabel metal1 4646 17136 4646 17136 0 _181_
rlabel metal1 6256 17238 6256 17238 0 _182_
rlabel metal2 6348 17102 6348 17102 0 _183_
rlabel metal2 7130 15776 7130 15776 0 _184_
rlabel metal1 6854 17136 6854 17136 0 _185_
rlabel metal1 6808 15130 6808 15130 0 _186_
rlabel metal1 6164 14518 6164 14518 0 _187_
rlabel metal2 5934 16116 5934 16116 0 _188_
rlabel metal1 5980 14246 5980 14246 0 _189_
rlabel metal1 5612 15538 5612 15538 0 _190_
rlabel metal1 6026 13192 6026 13192 0 _191_
rlabel metal2 4646 12444 4646 12444 0 _192_
rlabel metal1 4186 8874 4186 8874 0 _193_
rlabel metal1 3956 9010 3956 9010 0 _194_
rlabel metal1 3726 6630 3726 6630 0 _195_
rlabel viali 3626 6902 3626 6902 0 _196_
rlabel metal1 3358 6834 3358 6834 0 _197_
rlabel metal1 4554 5746 4554 5746 0 _198_
rlabel metal1 4370 5814 4370 5814 0 _199_
rlabel metal1 5198 5644 5198 5644 0 _200_
rlabel metal1 5382 5814 5382 5814 0 _201_
rlabel metal1 10166 3536 10166 3536 0 _202_
rlabel metal1 8694 6222 8694 6222 0 _203_
rlabel metal1 6118 7446 6118 7446 0 _204_
rlabel metal1 5566 8602 5566 8602 0 _205_
rlabel metal1 4968 11322 4968 11322 0 _206_
rlabel metal2 7222 13396 7222 13396 0 _207_
rlabel metal2 9706 14246 9706 14246 0 _208_
rlabel metal2 6486 11798 6486 11798 0 _209_
rlabel metal1 5704 12954 5704 12954 0 _210_
rlabel metal1 10534 15538 10534 15538 0 _211_
rlabel metal1 11546 14586 11546 14586 0 _212_
rlabel metal1 12604 16014 12604 16014 0 _213_
rlabel metal1 8694 16762 8694 16762 0 _214_
rlabel metal1 9798 17714 9798 17714 0 _215_
rlabel metal1 11224 17306 11224 17306 0 _216_
rlabel metal1 9798 15674 9798 15674 0 _217_
rlabel metal1 8188 14926 8188 14926 0 _218_
rlabel metal2 8418 9894 8418 9894 0 _219_
rlabel metal1 6762 6222 6762 6222 0 _220_
rlabel metal1 6762 5134 6762 5134 0 _221_
rlabel metal1 7544 3570 7544 3570 0 _222_
rlabel metal3 1970 17748 1970 17748 0 clk
rlabel metal1 6624 13838 6624 13838 0 clknet_0_clk
rlabel metal2 874 8160 874 8160 0 clknet_2_0__leaf_clk
rlabel metal2 12558 4046 12558 4046 0 clknet_2_1__leaf_clk
rlabel metal1 2346 14348 2346 14348 0 clknet_2_2__leaf_clk
rlabel metal1 10672 18258 10672 18258 0 clknet_2_3__leaf_clk
rlabel metal1 1364 3978 1364 3978 0 net1
rlabel metal1 15088 13974 15088 13974 0 net10
rlabel metal1 14766 13838 14766 13838 0 net11
rlabel metal1 14720 14450 14720 14450 0 net12
rlabel metal1 14628 13430 14628 13430 0 net13
rlabel metal1 11822 3978 11822 3978 0 net14
rlabel metal1 14536 782 14536 782 0 net15
rlabel metal2 2438 8670 2438 8670 0 net16
rlabel metal1 13156 3638 13156 3638 0 net17
rlabel metal2 2714 14620 2714 14620 0 net18
rlabel metal2 12558 17408 12558 17408 0 net19
rlabel metal2 17250 5100 17250 5100 0 net2
rlabel metal1 6341 14926 6341 14926 0 net20
rlabel via2 8050 12291 8050 12291 0 net21
rlabel metal1 5796 782 5796 782 0 net22
rlabel metal1 7498 1462 7498 1462 0 net23
rlabel metal1 10212 782 10212 782 0 net24
rlabel metal1 6486 2482 6486 2482 0 net25
rlabel metal1 6302 1938 6302 1938 0 net26
rlabel metal2 7222 2108 7222 2108 0 net27
rlabel metal1 6118 884 6118 884 0 net28
rlabel metal1 7820 918 7820 918 0 net29
rlabel metal1 17894 9520 17894 9520 0 net3
rlabel metal1 6762 2414 6762 2414 0 net30
rlabel metal1 5474 1428 5474 1428 0 net31
rlabel metal1 7820 986 7820 986 0 net32
rlabel metal1 8418 782 8418 782 0 net33
rlabel metal2 6578 1530 6578 1530 0 net34
rlabel metal1 7130 2482 7130 2482 0 net35
rlabel metal1 11730 1428 11730 1428 0 net36
rlabel metal2 7130 2244 7130 2244 0 net37
rlabel metal1 18860 12818 18860 12818 0 net38
rlabel metal3 590 1428 590 1428 0 net39
rlabel metal1 13570 5780 13570 5780 0 net4
rlabel metal2 3910 415 3910 415 0 net40
rlabel metal1 16192 18802 16192 18802 0 net41
rlabel metal2 19090 1547 19090 1547 0 net42
rlabel metal3 19328 1428 19328 1428 0 net43
rlabel metal1 19366 1394 19366 1394 0 net44
rlabel metal1 18124 18802 18124 18802 0 net45
rlabel metal1 15548 18802 15548 18802 0 net46
rlabel metal1 16008 8398 16008 8398 0 net47
rlabel metal3 590 18428 590 18428 0 net48
rlabel metal2 15502 500 15502 500 0 net49
rlabel metal1 13110 6154 13110 6154 0 net5
rlabel metal2 18078 500 18078 500 0 net50
rlabel metal1 3956 18938 3956 18938 0 net51
rlabel metal1 3128 4046 3128 4046 0 net52
rlabel metal1 1334 4046 1334 4046 0 net53
rlabel metal1 7958 2822 7958 2822 0 net54
rlabel metal1 8786 2074 8786 2074 0 net55
rlabel metal1 3726 3706 3726 3706 0 net56
rlabel metal1 10718 1530 10718 1530 0 net57
rlabel metal1 5474 15572 5474 15572 0 net58
rlabel metal1 5566 5678 5566 5678 0 net59
rlabel metal2 16606 3876 16606 3876 0 net6
rlabel metal1 2024 10574 2024 10574 0 net60
rlabel metal1 2162 6766 2162 6766 0 net61
rlabel metal2 3542 12954 3542 12954 0 net62
rlabel metal1 5060 17102 5060 17102 0 net63
rlabel metal2 1886 14892 1886 14892 0 net64
rlabel metal1 16376 4658 16376 4658 0 net65
rlabel metal1 7130 16218 7130 16218 0 net66
rlabel metal1 7728 1326 7728 1326 0 net67
rlabel metal1 13984 4998 13984 4998 0 net68
rlabel metal2 16514 11696 16514 11696 0 net69
rlabel metal2 13938 5610 13938 5610 0 net7
rlabel metal1 17204 14994 17204 14994 0 net70
rlabel metal1 13754 1870 13754 1870 0 net71
rlabel metal1 14398 2516 14398 2516 0 net72
rlabel metal2 8694 16014 8694 16014 0 net8
rlabel metal1 8050 8908 8050 8908 0 net9
rlabel metal1 2990 3570 2990 3570 0 res1_n
rlabel metal1 6118 5746 6118 5746 0 res2_n
rlabel metal3 406 4148 406 4148 0 rst_n
rlabel metal2 8878 4046 8878 4046 0 ts.o_res\[0\]
rlabel metal2 12098 14314 12098 14314 0 ts.o_res\[10\]
rlabel metal1 9384 16762 9384 16762 0 ts.o_res\[11\]
rlabel metal1 9154 18054 9154 18054 0 ts.o_res\[12\]
rlabel metal1 12926 13838 12926 13838 0 ts.o_res\[13\]
rlabel metal1 11040 15674 11040 15674 0 ts.o_res\[14\]
rlabel metal2 9246 15674 9246 15674 0 ts.o_res\[15\]
rlabel metal1 8326 9554 8326 9554 0 ts.o_res\[16\]
rlabel metal2 8786 8126 8786 8126 0 ts.o_res\[17\]
rlabel metal1 8694 7344 8694 7344 0 ts.o_res\[18\]
rlabel metal2 8142 8466 8142 8466 0 ts.o_res\[19\]
rlabel metal2 9154 8874 9154 8874 0 ts.o_res\[1\]
rlabel metal3 10235 12852 10235 12852 0 ts.o_res\[2\]
rlabel metal1 8970 9078 8970 9078 0 ts.o_res\[3\]
rlabel metal2 9338 10608 9338 10608 0 ts.o_res\[4\]
rlabel metal2 8142 13022 8142 13022 0 ts.o_res\[5\]
rlabel metal1 10028 13838 10028 13838 0 ts.o_res\[6\]
rlabel metal1 7268 11322 7268 11322 0 ts.o_res\[7\]
rlabel metal1 6394 12818 6394 12818 0 ts.o_res\[8\]
rlabel metal2 13386 14620 13386 14620 0 ts.o_res\[9\]
rlabel metal2 13754 7361 13754 7361 0 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal2 17526 4420 17526 4420 0 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal1 16974 4658 16974 4658 0 ts.ts_core.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal1 16974 8500 16974 8500 0 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal1 17342 7310 17342 7310 0 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal1 16376 9078 16376 9078 0 ts.ts_core.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal1 15870 4692 15870 4692 0 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal1 15134 3060 15134 3060 0 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal1 14076 5678 14076 5678 0 ts.ts_core.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal1 10212 3026 10212 3026 0 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal1 12926 2482 12926 2482 0 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal1 13248 6290 13248 6290 0 ts.ts_core.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal1 13616 4114 13616 4114 0 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal1 18216 11254 18216 11254 0 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal2 12374 5695 12374 5695 0 ts.ts_core.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal1 17158 8398 17158 8398 0 ts.ts_core.dac.vdac_single.en_pupd
rlabel metal1 15088 12818 15088 12818 0 ts.ts_core.dac_vout_ana_
rlabel metal1 11914 1428 11914 1428 0 ts.ts_core.dcdel_capnode_ana_
rlabel metal1 6565 1870 6565 1870 0 ts.ts_core.dcdel_out_n
rlabel metal1 14122 2006 14122 2006 0 ts.ts_core.i_precharge_n
rlabel metal4 12604 8500 12604 8500 0 ts.ts_core.o_tempdelay
rlabel metal1 6693 2074 6693 2074 0 ts.ts_core.tempdelay_async
rlabel metal2 11546 1836 11546 1836 0 ts.ts_core.tempdelay_sync1
rlabel metal1 13110 5678 13110 5678 0 ts.ts_ctrl.state\[0\]
rlabel metal1 13386 5542 13386 5542 0 ts.ts_ctrl.state\[1\]
rlabel metal1 7222 14892 7222 14892 0 ts.ts_ctrl.state\[2\]
rlabel metal1 10350 6970 10350 6970 0 ts.ts_ctrl.temp_ctr\[0\]
rlabel metal2 11546 14654 11546 14654 0 ts.ts_ctrl.temp_ctr\[10\]
rlabel metal1 6808 13974 6808 13974 0 ts.ts_ctrl.temp_ctr\[11\]
rlabel metal1 6808 13702 6808 13702 0 ts.ts_ctrl.temp_ctr\[12\]
rlabel metal1 11868 16966 11868 16966 0 ts.ts_ctrl.temp_ctr\[13\]
rlabel metal1 7866 15946 7866 15946 0 ts.ts_ctrl.temp_ctr\[14\]
rlabel metal1 6762 15028 6762 15028 0 ts.ts_ctrl.temp_ctr\[15\]
rlabel metal2 8786 9180 8786 9180 0 ts.ts_ctrl.temp_ctr\[16\]
rlabel metal1 7866 6154 7866 6154 0 ts.ts_ctrl.temp_ctr\[17\]
rlabel metal1 7682 5134 7682 5134 0 ts.ts_ctrl.temp_ctr\[18\]
rlabel metal1 7314 5644 7314 5644 0 ts.ts_ctrl.temp_ctr\[19\]
rlabel metal1 11086 7310 11086 7310 0 ts.ts_ctrl.temp_ctr\[1\]
rlabel metal1 2208 8330 2208 8330 0 ts.ts_ctrl.temp_ctr\[2\]
rlabel metal2 2622 8602 2622 8602 0 ts.ts_ctrl.temp_ctr\[3\]
rlabel metal1 5382 11322 5382 11322 0 ts.ts_ctrl.temp_ctr\[4\]
rlabel metal1 3496 12954 3496 12954 0 ts.ts_ctrl.temp_ctr\[5\]
rlabel metal1 5244 13294 5244 13294 0 ts.ts_ctrl.temp_ctr\[6\]
rlabel metal1 7130 11254 7130 11254 0 ts.ts_ctrl.temp_ctr\[7\]
rlabel metal1 7222 12614 7222 12614 0 ts.ts_ctrl.temp_ctr\[8\]
rlabel metal1 2346 14552 2346 14552 0 ts.ts_ctrl.temp_ctr\[9\]
rlabel metal2 19090 11351 19090 11351 0 ui_in[0]
rlabel metal1 18998 10574 18998 10574 0 ui_in[1]
rlabel metal1 18446 3502 18446 3502 0 ui_in[2]
rlabel metal1 18584 4046 18584 4046 0 ui_in[3]
rlabel metal1 19366 2482 19366 2482 0 ui_in[4]
rlabel metal1 19412 2958 19412 2958 0 ui_in[5]
rlabel metal1 8142 18870 8142 18870 0 ui_in[6]
rlabel metal1 18998 14348 18998 14348 0 ui_in[7]
rlabel metal1 19136 13838 19136 13838 0 uio_in[0]
rlabel metal1 19044 16014 19044 16014 0 uio_in[1]
rlabel metal2 18998 15487 18998 15487 0 uio_in[2]
rlabel metal1 19044 14858 19044 14858 0 uio_in[3]
rlabel metal2 10994 1557 10994 1557 0 uio_out[4]
rlabel metal2 15594 9333 15594 9333 0 uio_out[5]
rlabel metal2 12282 619 12282 619 0 uio_out[6]
rlabel metal2 15778 9775 15778 9775 0 uio_out[7]
rlabel metal1 8602 11254 8602 11254 0 uo_out[0]
rlabel metal1 12558 11118 12558 11118 0 uo_out[1]
rlabel via2 15134 11611 15134 11611 0 uo_out[2]
rlabel metal3 843 10948 843 10948 0 uo_out[3]
rlabel metal1 10074 18734 10074 18734 0 uo_out[4]
rlabel metal1 10304 12954 10304 12954 0 uo_out[5]
rlabel metal2 10810 15589 10810 15589 0 uo_out[6]
rlabel metal2 9062 16177 9062 16177 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
