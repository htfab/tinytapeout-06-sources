magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< nwell >>
rect -1199 -384 1199 384
<< pmos >>
rect -1003 -236 -803 164
rect -745 -236 -545 164
rect -487 -236 -287 164
rect -229 -236 -29 164
rect 29 -236 229 164
rect 287 -236 487 164
rect 545 -236 745 164
rect 803 -236 1003 164
<< pdiff >>
rect -1061 152 -1003 164
rect -1061 -224 -1049 152
rect -1015 -224 -1003 152
rect -1061 -236 -1003 -224
rect -803 152 -745 164
rect -803 -224 -791 152
rect -757 -224 -745 152
rect -803 -236 -745 -224
rect -545 152 -487 164
rect -545 -224 -533 152
rect -499 -224 -487 152
rect -545 -236 -487 -224
rect -287 152 -229 164
rect -287 -224 -275 152
rect -241 -224 -229 152
rect -287 -236 -229 -224
rect -29 152 29 164
rect -29 -224 -17 152
rect 17 -224 29 152
rect -29 -236 29 -224
rect 229 152 287 164
rect 229 -224 241 152
rect 275 -224 287 152
rect 229 -236 287 -224
rect 487 152 545 164
rect 487 -224 499 152
rect 533 -224 545 152
rect 487 -236 545 -224
rect 745 152 803 164
rect 745 -224 757 152
rect 791 -224 803 152
rect 745 -236 803 -224
rect 1003 152 1061 164
rect 1003 -224 1015 152
rect 1049 -224 1061 152
rect 1003 -236 1061 -224
<< pdiffc >>
rect -1049 -224 -1015 152
rect -791 -224 -757 152
rect -533 -224 -499 152
rect -275 -224 -241 152
rect -17 -224 17 152
rect 241 -224 275 152
rect 499 -224 533 152
rect 757 -224 791 152
rect 1015 -224 1049 152
<< nsubdiff >>
rect -1163 314 -1067 348
rect 1067 314 1163 348
rect -1163 -314 -1129 314
rect 1129 -314 1163 314
rect -1163 -348 1163 -314
<< nsubdiffcont >>
rect -1067 314 1067 348
<< poly >>
rect -1003 245 -803 261
rect -1003 211 -987 245
rect -819 211 -803 245
rect -1003 164 -803 211
rect -745 245 -545 261
rect -745 211 -729 245
rect -561 211 -545 245
rect -745 164 -545 211
rect -487 245 -287 261
rect -487 211 -471 245
rect -303 211 -287 245
rect -487 164 -287 211
rect -229 245 -29 261
rect -229 211 -213 245
rect -45 211 -29 245
rect -229 164 -29 211
rect 29 245 229 261
rect 29 211 45 245
rect 213 211 229 245
rect 29 164 229 211
rect 287 245 487 261
rect 287 211 303 245
rect 471 211 487 245
rect 287 164 487 211
rect 545 245 745 261
rect 545 211 561 245
rect 729 211 745 245
rect 545 164 745 211
rect 803 245 1003 261
rect 803 211 819 245
rect 987 211 1003 245
rect 803 164 1003 211
rect -1003 -262 -803 -236
rect -745 -262 -545 -236
rect -487 -262 -287 -236
rect -229 -262 -29 -236
rect 29 -262 229 -236
rect 287 -262 487 -236
rect 545 -262 745 -236
rect 803 -262 1003 -236
<< polycont >>
rect -987 211 -819 245
rect -729 211 -561 245
rect -471 211 -303 245
rect -213 211 -45 245
rect 45 211 213 245
rect 303 211 471 245
rect 561 211 729 245
rect 819 211 987 245
<< locali >>
rect -1163 -314 -1129 348
rect -1003 211 -987 245
rect -819 211 -803 245
rect -745 211 -729 245
rect -561 211 -545 245
rect -487 211 -471 245
rect -303 211 -287 245
rect -229 211 -213 245
rect -45 211 -29 245
rect 29 211 45 245
rect 213 211 229 245
rect 287 211 303 245
rect 471 211 487 245
rect 545 211 561 245
rect 729 211 745 245
rect 803 211 819 245
rect 987 211 1003 245
rect -1049 152 -1015 168
rect -1049 -240 -1015 -224
rect -791 152 -757 168
rect -791 -240 -757 -224
rect -533 152 -499 168
rect -533 -240 -499 -224
rect -275 152 -241 168
rect -275 -240 -241 -224
rect -17 152 17 168
rect -17 -240 17 -224
rect 241 152 275 168
rect 241 -240 275 -224
rect 499 152 533 168
rect 499 -240 533 -224
rect 757 152 791 168
rect 757 -240 791 -224
rect 1015 152 1049 168
rect 1015 -240 1049 -224
rect 1129 -314 1163 348
rect -1163 -348 1163 -314
<< viali >>
rect -1129 314 -1067 348
rect -1067 314 1067 348
rect 1067 314 1129 348
rect -987 211 -819 245
rect -729 211 -561 245
rect -471 211 -303 245
rect -213 211 -45 245
rect 45 211 213 245
rect 303 211 471 245
rect 561 211 729 245
rect 819 211 987 245
rect -1049 -224 -1015 152
rect -791 -224 -757 152
rect -533 -224 -499 152
rect -275 -224 -241 152
rect -17 -224 17 152
rect 241 -224 275 152
rect 499 -224 533 152
rect 757 -224 791 152
rect 1015 -224 1049 152
<< metal1 >>
rect -1141 348 1141 354
rect -1141 314 -1129 348
rect 1129 314 1141 348
rect -1141 308 1141 314
rect -999 245 -807 251
rect -999 211 -987 245
rect -819 211 -807 245
rect -999 205 -807 211
rect -741 245 -549 251
rect -741 211 -729 245
rect -561 211 -549 245
rect -741 205 -549 211
rect -483 245 -291 251
rect -483 211 -471 245
rect -303 211 -291 245
rect -483 205 -291 211
rect -225 245 -33 251
rect -225 211 -213 245
rect -45 211 -33 245
rect -225 205 -33 211
rect 33 245 225 251
rect 33 211 45 245
rect 213 211 225 245
rect 33 205 225 211
rect 291 245 483 251
rect 291 211 303 245
rect 471 211 483 245
rect 291 205 483 211
rect 549 245 741 251
rect 549 211 561 245
rect 729 211 741 245
rect 549 205 741 211
rect 807 245 999 251
rect 807 211 819 245
rect 987 211 999 245
rect 807 205 999 211
rect -1055 152 -1009 164
rect -1055 -224 -1049 152
rect -1015 -224 -1009 152
rect -1055 -236 -1009 -224
rect -797 152 -751 164
rect -797 -224 -791 152
rect -757 -224 -751 152
rect -797 -236 -751 -224
rect -539 152 -493 164
rect -539 -224 -533 152
rect -499 -224 -493 152
rect -539 -236 -493 -224
rect -281 152 -235 164
rect -281 -224 -275 152
rect -241 -224 -235 152
rect -281 -236 -235 -224
rect -23 152 23 164
rect -23 -224 -17 152
rect 17 -224 23 152
rect -23 -236 23 -224
rect 235 152 281 164
rect 235 -224 241 152
rect 275 -224 281 152
rect 235 -236 281 -224
rect 493 152 539 164
rect 493 -224 499 152
rect 533 -224 539 152
rect 493 -236 539 -224
rect 751 152 797 164
rect 751 -224 757 152
rect 791 -224 797 152
rect 751 -236 797 -224
rect 1009 152 1055 164
rect 1009 -224 1015 152
rect 1049 -224 1055 152
rect 1009 -236 1055 -224
<< properties >>
string FIXED_BBOX -1146 -331 1146 331
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
