magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -2231 -719 2231 719
<< nmos >>
rect -2035 109 -1835 509
rect -1777 109 -1577 509
rect -1519 109 -1319 509
rect -1261 109 -1061 509
rect -1003 109 -803 509
rect -745 109 -545 509
rect -487 109 -287 509
rect -229 109 -29 509
rect 29 109 229 509
rect 287 109 487 509
rect 545 109 745 509
rect 803 109 1003 509
rect 1061 109 1261 509
rect 1319 109 1519 509
rect 1577 109 1777 509
rect 1835 109 2035 509
rect -2035 -509 -1835 -109
rect -1777 -509 -1577 -109
rect -1519 -509 -1319 -109
rect -1261 -509 -1061 -109
rect -1003 -509 -803 -109
rect -745 -509 -545 -109
rect -487 -509 -287 -109
rect -229 -509 -29 -109
rect 29 -509 229 -109
rect 287 -509 487 -109
rect 545 -509 745 -109
rect 803 -509 1003 -109
rect 1061 -509 1261 -109
rect 1319 -509 1519 -109
rect 1577 -509 1777 -109
rect 1835 -509 2035 -109
<< ndiff >>
rect -2093 497 -2035 509
rect -2093 121 -2081 497
rect -2047 121 -2035 497
rect -2093 109 -2035 121
rect -1835 497 -1777 509
rect -1835 121 -1823 497
rect -1789 121 -1777 497
rect -1835 109 -1777 121
rect -1577 497 -1519 509
rect -1577 121 -1565 497
rect -1531 121 -1519 497
rect -1577 109 -1519 121
rect -1319 497 -1261 509
rect -1319 121 -1307 497
rect -1273 121 -1261 497
rect -1319 109 -1261 121
rect -1061 497 -1003 509
rect -1061 121 -1049 497
rect -1015 121 -1003 497
rect -1061 109 -1003 121
rect -803 497 -745 509
rect -803 121 -791 497
rect -757 121 -745 497
rect -803 109 -745 121
rect -545 497 -487 509
rect -545 121 -533 497
rect -499 121 -487 497
rect -545 109 -487 121
rect -287 497 -229 509
rect -287 121 -275 497
rect -241 121 -229 497
rect -287 109 -229 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 229 497 287 509
rect 229 121 241 497
rect 275 121 287 497
rect 229 109 287 121
rect 487 497 545 509
rect 487 121 499 497
rect 533 121 545 497
rect 487 109 545 121
rect 745 497 803 509
rect 745 121 757 497
rect 791 121 803 497
rect 745 109 803 121
rect 1003 497 1061 509
rect 1003 121 1015 497
rect 1049 121 1061 497
rect 1003 109 1061 121
rect 1261 497 1319 509
rect 1261 121 1273 497
rect 1307 121 1319 497
rect 1261 109 1319 121
rect 1519 497 1577 509
rect 1519 121 1531 497
rect 1565 121 1577 497
rect 1519 109 1577 121
rect 1777 497 1835 509
rect 1777 121 1789 497
rect 1823 121 1835 497
rect 1777 109 1835 121
rect 2035 497 2093 509
rect 2035 121 2047 497
rect 2081 121 2093 497
rect 2035 109 2093 121
rect -2093 -121 -2035 -109
rect -2093 -497 -2081 -121
rect -2047 -497 -2035 -121
rect -2093 -509 -2035 -497
rect -1835 -121 -1777 -109
rect -1835 -497 -1823 -121
rect -1789 -497 -1777 -121
rect -1835 -509 -1777 -497
rect -1577 -121 -1519 -109
rect -1577 -497 -1565 -121
rect -1531 -497 -1519 -121
rect -1577 -509 -1519 -497
rect -1319 -121 -1261 -109
rect -1319 -497 -1307 -121
rect -1273 -497 -1261 -121
rect -1319 -509 -1261 -497
rect -1061 -121 -1003 -109
rect -1061 -497 -1049 -121
rect -1015 -497 -1003 -121
rect -1061 -509 -1003 -497
rect -803 -121 -745 -109
rect -803 -497 -791 -121
rect -757 -497 -745 -121
rect -803 -509 -745 -497
rect -545 -121 -487 -109
rect -545 -497 -533 -121
rect -499 -497 -487 -121
rect -545 -509 -487 -497
rect -287 -121 -229 -109
rect -287 -497 -275 -121
rect -241 -497 -229 -121
rect -287 -509 -229 -497
rect -29 -121 29 -109
rect -29 -497 -17 -121
rect 17 -497 29 -121
rect -29 -509 29 -497
rect 229 -121 287 -109
rect 229 -497 241 -121
rect 275 -497 287 -121
rect 229 -509 287 -497
rect 487 -121 545 -109
rect 487 -497 499 -121
rect 533 -497 545 -121
rect 487 -509 545 -497
rect 745 -121 803 -109
rect 745 -497 757 -121
rect 791 -497 803 -121
rect 745 -509 803 -497
rect 1003 -121 1061 -109
rect 1003 -497 1015 -121
rect 1049 -497 1061 -121
rect 1003 -509 1061 -497
rect 1261 -121 1319 -109
rect 1261 -497 1273 -121
rect 1307 -497 1319 -121
rect 1261 -509 1319 -497
rect 1519 -121 1577 -109
rect 1519 -497 1531 -121
rect 1565 -497 1577 -121
rect 1519 -509 1577 -497
rect 1777 -121 1835 -109
rect 1777 -497 1789 -121
rect 1823 -497 1835 -121
rect 1777 -509 1835 -497
rect 2035 -121 2093 -109
rect 2035 -497 2047 -121
rect 2081 -497 2093 -121
rect 2035 -509 2093 -497
<< ndiffc >>
rect -2081 121 -2047 497
rect -1823 121 -1789 497
rect -1565 121 -1531 497
rect -1307 121 -1273 497
rect -1049 121 -1015 497
rect -791 121 -757 497
rect -533 121 -499 497
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect 499 121 533 497
rect 757 121 791 497
rect 1015 121 1049 497
rect 1273 121 1307 497
rect 1531 121 1565 497
rect 1789 121 1823 497
rect 2047 121 2081 497
rect -2081 -497 -2047 -121
rect -1823 -497 -1789 -121
rect -1565 -497 -1531 -121
rect -1307 -497 -1273 -121
rect -1049 -497 -1015 -121
rect -791 -497 -757 -121
rect -533 -497 -499 -121
rect -275 -497 -241 -121
rect -17 -497 17 -121
rect 241 -497 275 -121
rect 499 -497 533 -121
rect 757 -497 791 -121
rect 1015 -497 1049 -121
rect 1273 -497 1307 -121
rect 1531 -497 1565 -121
rect 1789 -497 1823 -121
rect 2047 -497 2081 -121
<< psubdiff >>
rect -2195 649 2195 683
rect -2195 587 -2161 649
rect 2161 587 2195 649
rect -2195 -649 -2161 -587
rect 2161 -649 2195 -587
rect -2195 -683 -2099 -649
rect 2099 -683 2195 -649
<< psubdiffcont >>
rect -2195 -587 -2161 587
rect 2161 -587 2195 587
rect -2099 -683 2099 -649
<< poly >>
rect -2035 581 -1835 597
rect -2035 547 -2019 581
rect -1851 547 -1835 581
rect -2035 509 -1835 547
rect -1777 581 -1577 597
rect -1777 547 -1761 581
rect -1593 547 -1577 581
rect -1777 509 -1577 547
rect -1519 581 -1319 597
rect -1519 547 -1503 581
rect -1335 547 -1319 581
rect -1519 509 -1319 547
rect -1261 581 -1061 597
rect -1261 547 -1245 581
rect -1077 547 -1061 581
rect -1261 509 -1061 547
rect -1003 581 -803 597
rect -1003 547 -987 581
rect -819 547 -803 581
rect -1003 509 -803 547
rect -745 581 -545 597
rect -745 547 -729 581
rect -561 547 -545 581
rect -745 509 -545 547
rect -487 581 -287 597
rect -487 547 -471 581
rect -303 547 -287 581
rect -487 509 -287 547
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 509 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 509 229 547
rect 287 581 487 597
rect 287 547 303 581
rect 471 547 487 581
rect 287 509 487 547
rect 545 581 745 597
rect 545 547 561 581
rect 729 547 745 581
rect 545 509 745 547
rect 803 581 1003 597
rect 803 547 819 581
rect 987 547 1003 581
rect 803 509 1003 547
rect 1061 581 1261 597
rect 1061 547 1077 581
rect 1245 547 1261 581
rect 1061 509 1261 547
rect 1319 581 1519 597
rect 1319 547 1335 581
rect 1503 547 1519 581
rect 1319 509 1519 547
rect 1577 581 1777 597
rect 1577 547 1593 581
rect 1761 547 1777 581
rect 1577 509 1777 547
rect 1835 581 2035 597
rect 1835 547 1851 581
rect 2019 547 2035 581
rect 1835 509 2035 547
rect -2035 71 -1835 109
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 109
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 109
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 109
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 109
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 109
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 109
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 109
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -109 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -109 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -109 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -109 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -109 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -109 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -109 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -109 2035 -71
rect -2035 -547 -1835 -509
rect -2035 -581 -2019 -547
rect -1851 -581 -1835 -547
rect -2035 -597 -1835 -581
rect -1777 -547 -1577 -509
rect -1777 -581 -1761 -547
rect -1593 -581 -1577 -547
rect -1777 -597 -1577 -581
rect -1519 -547 -1319 -509
rect -1519 -581 -1503 -547
rect -1335 -581 -1319 -547
rect -1519 -597 -1319 -581
rect -1261 -547 -1061 -509
rect -1261 -581 -1245 -547
rect -1077 -581 -1061 -547
rect -1261 -597 -1061 -581
rect -1003 -547 -803 -509
rect -1003 -581 -987 -547
rect -819 -581 -803 -547
rect -1003 -597 -803 -581
rect -745 -547 -545 -509
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -745 -597 -545 -581
rect -487 -547 -287 -509
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -487 -597 -287 -581
rect -229 -547 -29 -509
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -509
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
rect 287 -547 487 -509
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 287 -597 487 -581
rect 545 -547 745 -509
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 545 -597 745 -581
rect 803 -547 1003 -509
rect 803 -581 819 -547
rect 987 -581 1003 -547
rect 803 -597 1003 -581
rect 1061 -547 1261 -509
rect 1061 -581 1077 -547
rect 1245 -581 1261 -547
rect 1061 -597 1261 -581
rect 1319 -547 1519 -509
rect 1319 -581 1335 -547
rect 1503 -581 1519 -547
rect 1319 -597 1519 -581
rect 1577 -547 1777 -509
rect 1577 -581 1593 -547
rect 1761 -581 1777 -547
rect 1577 -597 1777 -581
rect 1835 -547 2035 -509
rect 1835 -581 1851 -547
rect 2019 -581 2035 -547
rect 1835 -597 2035 -581
<< polycont >>
rect -2019 547 -1851 581
rect -1761 547 -1593 581
rect -1503 547 -1335 581
rect -1245 547 -1077 581
rect -987 547 -819 581
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect 819 547 987 581
rect 1077 547 1245 581
rect 1335 547 1503 581
rect 1593 547 1761 581
rect 1851 547 2019 581
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect -2019 -581 -1851 -547
rect -1761 -581 -1593 -547
rect -1503 -581 -1335 -547
rect -1245 -581 -1077 -547
rect -987 -581 -819 -547
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
rect 819 -581 987 -547
rect 1077 -581 1245 -547
rect 1335 -581 1503 -547
rect 1593 -581 1761 -547
rect 1851 -581 2019 -547
<< locali >>
rect -2195 587 -2161 683
rect 2161 587 2195 683
rect -2035 547 -2019 581
rect -1851 547 -1835 581
rect -1777 547 -1761 581
rect -1593 547 -1577 581
rect -1519 547 -1503 581
rect -1335 547 -1319 581
rect -1261 547 -1245 581
rect -1077 547 -1061 581
rect -1003 547 -987 581
rect -819 547 -803 581
rect -745 547 -729 581
rect -561 547 -545 581
rect -487 547 -471 581
rect -303 547 -287 581
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect 287 547 303 581
rect 471 547 487 581
rect 545 547 561 581
rect 729 547 745 581
rect 803 547 819 581
rect 987 547 1003 581
rect 1061 547 1077 581
rect 1245 547 1261 581
rect 1319 547 1335 581
rect 1503 547 1519 581
rect 1577 547 1593 581
rect 1761 547 1777 581
rect 1835 547 1851 581
rect 2019 547 2035 581
rect -2081 497 -2047 513
rect -2081 105 -2047 121
rect -1823 497 -1789 513
rect -1823 105 -1789 121
rect -1565 497 -1531 513
rect -1565 105 -1531 121
rect -1307 497 -1273 513
rect -1307 105 -1273 121
rect -1049 497 -1015 513
rect -1049 105 -1015 121
rect -791 497 -757 513
rect -791 105 -757 121
rect -533 497 -499 513
rect -533 105 -499 121
rect -275 497 -241 513
rect -275 105 -241 121
rect -17 497 17 513
rect -17 105 17 121
rect 241 497 275 513
rect 241 105 275 121
rect 499 497 533 513
rect 499 105 533 121
rect 757 497 791 513
rect 757 105 791 121
rect 1015 497 1049 513
rect 1015 105 1049 121
rect 1273 497 1307 513
rect 1273 105 1307 121
rect 1531 497 1565 513
rect 1531 105 1565 121
rect 1789 497 1823 513
rect 1789 105 1823 121
rect 2047 497 2081 513
rect 2047 105 2081 121
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect -2081 -121 -2047 -105
rect -2081 -513 -2047 -497
rect -1823 -121 -1789 -105
rect -1823 -513 -1789 -497
rect -1565 -121 -1531 -105
rect -1565 -513 -1531 -497
rect -1307 -121 -1273 -105
rect -1307 -513 -1273 -497
rect -1049 -121 -1015 -105
rect -1049 -513 -1015 -497
rect -791 -121 -757 -105
rect -791 -513 -757 -497
rect -533 -121 -499 -105
rect -533 -513 -499 -497
rect -275 -121 -241 -105
rect -275 -513 -241 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 241 -121 275 -105
rect 241 -513 275 -497
rect 499 -121 533 -105
rect 499 -513 533 -497
rect 757 -121 791 -105
rect 757 -513 791 -497
rect 1015 -121 1049 -105
rect 1015 -513 1049 -497
rect 1273 -121 1307 -105
rect 1273 -513 1307 -497
rect 1531 -121 1565 -105
rect 1531 -513 1565 -497
rect 1789 -121 1823 -105
rect 1789 -513 1823 -497
rect 2047 -121 2081 -105
rect 2047 -513 2081 -497
rect -2035 -581 -2019 -547
rect -1851 -581 -1835 -547
rect -1777 -581 -1761 -547
rect -1593 -581 -1577 -547
rect -1519 -581 -1503 -547
rect -1335 -581 -1319 -547
rect -1261 -581 -1245 -547
rect -1077 -581 -1061 -547
rect -1003 -581 -987 -547
rect -819 -581 -803 -547
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 803 -581 819 -547
rect 987 -581 1003 -547
rect 1061 -581 1077 -547
rect 1245 -581 1261 -547
rect 1319 -581 1335 -547
rect 1503 -581 1519 -547
rect 1577 -581 1593 -547
rect 1761 -581 1777 -547
rect 1835 -581 1851 -547
rect 2019 -581 2035 -547
rect -2195 -683 -2099 -649
rect 2099 -683 2195 -649
<< viali >>
rect -2161 649 2161 683
rect -2019 547 -1851 581
rect -1761 547 -1593 581
rect -1503 547 -1335 581
rect -1245 547 -1077 581
rect -987 547 -819 581
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect 819 547 987 581
rect 1077 547 1245 581
rect 1335 547 1503 581
rect 1593 547 1761 581
rect 1851 547 2019 581
rect -2081 330 -2047 480
rect -1823 138 -1789 288
rect -1565 330 -1531 480
rect -1307 138 -1273 288
rect -1049 330 -1015 480
rect -791 138 -757 288
rect -533 330 -499 480
rect -275 138 -241 288
rect -17 330 17 480
rect 241 138 275 288
rect 499 330 533 480
rect 757 138 791 288
rect 1015 330 1049 480
rect 1273 138 1307 288
rect 1531 330 1565 480
rect 1789 138 1823 288
rect 2047 330 2081 480
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect -2195 -587 -2161 -130
rect -2081 -288 -2047 -138
rect -1823 -480 -1789 -330
rect -1565 -288 -1531 -138
rect -1307 -480 -1273 -330
rect -1049 -288 -1015 -138
rect -791 -480 -757 -330
rect -533 -288 -499 -138
rect -275 -480 -241 -330
rect -17 -288 17 -138
rect 241 -480 275 -330
rect 499 -288 533 -138
rect 757 -480 791 -330
rect 1015 -288 1049 -138
rect 1273 -480 1307 -330
rect 1531 -288 1565 -138
rect 1789 -480 1823 -330
rect 2047 -288 2081 -138
rect -2019 -581 -1851 -547
rect -1761 -581 -1593 -547
rect -1503 -581 -1335 -547
rect -1245 -581 -1077 -547
rect -987 -581 -819 -547
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
rect 819 -581 987 -547
rect 1077 -581 1245 -547
rect 1335 -581 1503 -547
rect 1593 -581 1761 -547
rect 1851 -581 2019 -547
rect -2195 -649 -2161 -587
rect 2161 -587 2195 -130
rect 2161 -649 2195 -587
<< metal1 >>
rect -2173 683 2173 689
rect -2173 649 -2161 683
rect 2161 649 2173 683
rect -2173 643 2173 649
rect -2031 581 -1839 587
rect -2031 547 -2019 581
rect -1851 547 -1839 581
rect -2031 541 -1839 547
rect -1773 581 -1581 587
rect -1773 547 -1761 581
rect -1593 547 -1581 581
rect -1773 541 -1581 547
rect -1515 581 -1323 587
rect -1515 547 -1503 581
rect -1335 547 -1323 581
rect -1515 541 -1323 547
rect -1257 581 -1065 587
rect -1257 547 -1245 581
rect -1077 547 -1065 581
rect -1257 541 -1065 547
rect -999 581 -807 587
rect -999 547 -987 581
rect -819 547 -807 581
rect -999 541 -807 547
rect -741 581 -549 587
rect -741 547 -729 581
rect -561 547 -549 581
rect -741 541 -549 547
rect -483 581 -291 587
rect -483 547 -471 581
rect -303 547 -291 581
rect -483 541 -291 547
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect 291 581 483 587
rect 291 547 303 581
rect 471 547 483 581
rect 291 541 483 547
rect 549 581 741 587
rect 549 547 561 581
rect 729 547 741 581
rect 549 541 741 547
rect 807 581 999 587
rect 807 547 819 581
rect 987 547 999 581
rect 807 541 999 547
rect 1065 581 1257 587
rect 1065 547 1077 581
rect 1245 547 1257 581
rect 1065 541 1257 547
rect 1323 581 1515 587
rect 1323 547 1335 581
rect 1503 547 1515 581
rect 1323 541 1515 547
rect 1581 581 1773 587
rect 1581 547 1593 581
rect 1761 547 1773 581
rect 1581 541 1773 547
rect 1839 581 2031 587
rect 1839 547 1851 581
rect 2019 547 2031 581
rect 1839 541 2031 547
rect -2087 480 -2041 492
rect -2087 330 -2081 480
rect -2047 330 -2041 480
rect -2087 318 -2041 330
rect -1571 480 -1525 492
rect -1571 330 -1565 480
rect -1531 330 -1525 480
rect -1571 318 -1525 330
rect -1055 480 -1009 492
rect -1055 330 -1049 480
rect -1015 330 -1009 480
rect -1055 318 -1009 330
rect -539 480 -493 492
rect -539 330 -533 480
rect -499 330 -493 480
rect -539 318 -493 330
rect -23 480 23 492
rect -23 330 -17 480
rect 17 330 23 480
rect -23 318 23 330
rect 493 480 539 492
rect 493 330 499 480
rect 533 330 539 480
rect 493 318 539 330
rect 1009 480 1055 492
rect 1009 330 1015 480
rect 1049 330 1055 480
rect 1009 318 1055 330
rect 1525 480 1571 492
rect 1525 330 1531 480
rect 1565 330 1571 480
rect 1525 318 1571 330
rect 2041 480 2087 492
rect 2041 330 2047 480
rect 2081 330 2087 480
rect 2041 318 2087 330
rect -1829 288 -1783 300
rect -1829 138 -1823 288
rect -1789 138 -1783 288
rect -1829 126 -1783 138
rect -1313 288 -1267 300
rect -1313 138 -1307 288
rect -1273 138 -1267 288
rect -1313 126 -1267 138
rect -797 288 -751 300
rect -797 138 -791 288
rect -757 138 -751 288
rect -797 126 -751 138
rect -281 288 -235 300
rect -281 138 -275 288
rect -241 138 -235 288
rect -281 126 -235 138
rect 235 288 281 300
rect 235 138 241 288
rect 275 138 281 288
rect 235 126 281 138
rect 751 288 797 300
rect 751 138 757 288
rect 791 138 797 288
rect 751 126 797 138
rect 1267 288 1313 300
rect 1267 138 1273 288
rect 1307 138 1313 288
rect 1267 126 1313 138
rect 1783 288 1829 300
rect 1783 138 1789 288
rect 1823 138 1829 288
rect 1783 126 1829 138
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect -2201 -130 -2155 -118
rect -2201 -649 -2195 -130
rect -2161 -649 -2155 -130
rect -2087 -138 -2041 -126
rect -2087 -288 -2081 -138
rect -2047 -288 -2041 -138
rect -2087 -300 -2041 -288
rect -1571 -138 -1525 -126
rect -1571 -288 -1565 -138
rect -1531 -288 -1525 -138
rect -1571 -300 -1525 -288
rect -1055 -138 -1009 -126
rect -1055 -288 -1049 -138
rect -1015 -288 -1009 -138
rect -1055 -300 -1009 -288
rect -539 -138 -493 -126
rect -539 -288 -533 -138
rect -499 -288 -493 -138
rect -539 -300 -493 -288
rect -23 -138 23 -126
rect -23 -288 -17 -138
rect 17 -288 23 -138
rect -23 -300 23 -288
rect 493 -138 539 -126
rect 493 -288 499 -138
rect 533 -288 539 -138
rect 493 -300 539 -288
rect 1009 -138 1055 -126
rect 1009 -288 1015 -138
rect 1049 -288 1055 -138
rect 1009 -300 1055 -288
rect 1525 -138 1571 -126
rect 1525 -288 1531 -138
rect 1565 -288 1571 -138
rect 1525 -300 1571 -288
rect 2041 -138 2087 -126
rect 2041 -288 2047 -138
rect 2081 -288 2087 -138
rect 2041 -300 2087 -288
rect 2155 -130 2201 -118
rect -1829 -330 -1783 -318
rect -1829 -480 -1823 -330
rect -1789 -480 -1783 -330
rect -1829 -492 -1783 -480
rect -1313 -330 -1267 -318
rect -1313 -480 -1307 -330
rect -1273 -480 -1267 -330
rect -1313 -492 -1267 -480
rect -797 -330 -751 -318
rect -797 -480 -791 -330
rect -757 -480 -751 -330
rect -797 -492 -751 -480
rect -281 -330 -235 -318
rect -281 -480 -275 -330
rect -241 -480 -235 -330
rect -281 -492 -235 -480
rect 235 -330 281 -318
rect 235 -480 241 -330
rect 275 -480 281 -330
rect 235 -492 281 -480
rect 751 -330 797 -318
rect 751 -480 757 -330
rect 791 -480 797 -330
rect 751 -492 797 -480
rect 1267 -330 1313 -318
rect 1267 -480 1273 -330
rect 1307 -480 1313 -330
rect 1267 -492 1313 -480
rect 1783 -330 1829 -318
rect 1783 -480 1789 -330
rect 1823 -480 1829 -330
rect 1783 -492 1829 -480
rect -2031 -547 -1839 -541
rect -2031 -581 -2019 -547
rect -1851 -581 -1839 -547
rect -2031 -587 -1839 -581
rect -1773 -547 -1581 -541
rect -1773 -581 -1761 -547
rect -1593 -581 -1581 -547
rect -1773 -587 -1581 -581
rect -1515 -547 -1323 -541
rect -1515 -581 -1503 -547
rect -1335 -581 -1323 -547
rect -1515 -587 -1323 -581
rect -1257 -547 -1065 -541
rect -1257 -581 -1245 -547
rect -1077 -581 -1065 -547
rect -1257 -587 -1065 -581
rect -999 -547 -807 -541
rect -999 -581 -987 -547
rect -819 -581 -807 -547
rect -999 -587 -807 -581
rect -741 -547 -549 -541
rect -741 -581 -729 -547
rect -561 -581 -549 -547
rect -741 -587 -549 -581
rect -483 -547 -291 -541
rect -483 -581 -471 -547
rect -303 -581 -291 -547
rect -483 -587 -291 -581
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
rect 291 -547 483 -541
rect 291 -581 303 -547
rect 471 -581 483 -547
rect 291 -587 483 -581
rect 549 -547 741 -541
rect 549 -581 561 -547
rect 729 -581 741 -547
rect 549 -587 741 -581
rect 807 -547 999 -541
rect 807 -581 819 -547
rect 987 -581 999 -547
rect 807 -587 999 -581
rect 1065 -547 1257 -541
rect 1065 -581 1077 -547
rect 1245 -581 1257 -547
rect 1065 -587 1257 -581
rect 1323 -547 1515 -541
rect 1323 -581 1335 -547
rect 1503 -581 1515 -547
rect 1323 -587 1515 -581
rect 1581 -547 1773 -541
rect 1581 -581 1593 -547
rect 1761 -581 1773 -547
rect 1581 -587 1773 -581
rect 1839 -547 2031 -541
rect 1839 -581 1851 -547
rect 2019 -581 2031 -547
rect 1839 -587 2031 -581
rect -2201 -661 -2155 -649
rect 2155 -649 2161 -130
rect 2195 -649 2201 -130
rect 2155 -661 2201 -649
<< properties >>
string FIXED_BBOX -2178 -666 2178 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
