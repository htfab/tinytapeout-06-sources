magic
tech sky130A
magscale 1 2
timestamp 1713055061
<< pwell >>
rect -2102 -657 2102 657
<< nmos >>
rect -1906 109 -1706 509
rect -1648 109 -1448 509
rect -1390 109 -1190 509
rect -1132 109 -932 509
rect -874 109 -674 509
rect -616 109 -416 509
rect -358 109 -158 509
rect -100 109 100 509
rect 158 109 358 509
rect 416 109 616 509
rect 674 109 874 509
rect 932 109 1132 509
rect 1190 109 1390 509
rect 1448 109 1648 509
rect 1706 109 1906 509
rect -1906 -447 -1706 -47
rect -1648 -447 -1448 -47
rect -1390 -447 -1190 -47
rect -1132 -447 -932 -47
rect -874 -447 -674 -47
rect -616 -447 -416 -47
rect -358 -447 -158 -47
rect -100 -447 100 -47
rect 158 -447 358 -47
rect 416 -447 616 -47
rect 674 -447 874 -47
rect 932 -447 1132 -47
rect 1190 -447 1390 -47
rect 1448 -447 1648 -47
rect 1706 -447 1906 -47
<< ndiff >>
rect -1964 497 -1906 509
rect -1964 121 -1952 497
rect -1918 121 -1906 497
rect -1964 109 -1906 121
rect -1706 497 -1648 509
rect -1706 121 -1694 497
rect -1660 121 -1648 497
rect -1706 109 -1648 121
rect -1448 497 -1390 509
rect -1448 121 -1436 497
rect -1402 121 -1390 497
rect -1448 109 -1390 121
rect -1190 497 -1132 509
rect -1190 121 -1178 497
rect -1144 121 -1132 497
rect -1190 109 -1132 121
rect -932 497 -874 509
rect -932 121 -920 497
rect -886 121 -874 497
rect -932 109 -874 121
rect -674 497 -616 509
rect -674 121 -662 497
rect -628 121 -616 497
rect -674 109 -616 121
rect -416 497 -358 509
rect -416 121 -404 497
rect -370 121 -358 497
rect -416 109 -358 121
rect -158 497 -100 509
rect -158 121 -146 497
rect -112 121 -100 497
rect -158 109 -100 121
rect 100 497 158 509
rect 100 121 112 497
rect 146 121 158 497
rect 100 109 158 121
rect 358 497 416 509
rect 358 121 370 497
rect 404 121 416 497
rect 358 109 416 121
rect 616 497 674 509
rect 616 121 628 497
rect 662 121 674 497
rect 616 109 674 121
rect 874 497 932 509
rect 874 121 886 497
rect 920 121 932 497
rect 874 109 932 121
rect 1132 497 1190 509
rect 1132 121 1144 497
rect 1178 121 1190 497
rect 1132 109 1190 121
rect 1390 497 1448 509
rect 1390 121 1402 497
rect 1436 121 1448 497
rect 1390 109 1448 121
rect 1648 497 1706 509
rect 1648 121 1660 497
rect 1694 121 1706 497
rect 1648 109 1706 121
rect 1906 497 1964 509
rect 1906 121 1918 497
rect 1952 121 1964 497
rect 1906 109 1964 121
rect -1964 -59 -1906 -47
rect -1964 -435 -1952 -59
rect -1918 -435 -1906 -59
rect -1964 -447 -1906 -435
rect -1706 -59 -1648 -47
rect -1706 -435 -1694 -59
rect -1660 -435 -1648 -59
rect -1706 -447 -1648 -435
rect -1448 -59 -1390 -47
rect -1448 -435 -1436 -59
rect -1402 -435 -1390 -59
rect -1448 -447 -1390 -435
rect -1190 -59 -1132 -47
rect -1190 -435 -1178 -59
rect -1144 -435 -1132 -59
rect -1190 -447 -1132 -435
rect -932 -59 -874 -47
rect -932 -435 -920 -59
rect -886 -435 -874 -59
rect -932 -447 -874 -435
rect -674 -59 -616 -47
rect -674 -435 -662 -59
rect -628 -435 -616 -59
rect -674 -447 -616 -435
rect -416 -59 -358 -47
rect -416 -435 -404 -59
rect -370 -435 -358 -59
rect -416 -447 -358 -435
rect -158 -59 -100 -47
rect -158 -435 -146 -59
rect -112 -435 -100 -59
rect -158 -447 -100 -435
rect 100 -59 158 -47
rect 100 -435 112 -59
rect 146 -435 158 -59
rect 100 -447 158 -435
rect 358 -59 416 -47
rect 358 -435 370 -59
rect 404 -435 416 -59
rect 358 -447 416 -435
rect 616 -59 674 -47
rect 616 -435 628 -59
rect 662 -435 674 -59
rect 616 -447 674 -435
rect 874 -59 932 -47
rect 874 -435 886 -59
rect 920 -435 932 -59
rect 874 -447 932 -435
rect 1132 -59 1190 -47
rect 1132 -435 1144 -59
rect 1178 -435 1190 -59
rect 1132 -447 1190 -435
rect 1390 -59 1448 -47
rect 1390 -435 1402 -59
rect 1436 -435 1448 -59
rect 1390 -447 1448 -435
rect 1648 -59 1706 -47
rect 1648 -435 1660 -59
rect 1694 -435 1706 -59
rect 1648 -447 1706 -435
rect 1906 -59 1964 -47
rect 1906 -435 1918 -59
rect 1952 -435 1964 -59
rect 1906 -447 1964 -435
<< ndiffc >>
rect -1952 121 -1918 497
rect -1694 121 -1660 497
rect -1436 121 -1402 497
rect -1178 121 -1144 497
rect -920 121 -886 497
rect -662 121 -628 497
rect -404 121 -370 497
rect -146 121 -112 497
rect 112 121 146 497
rect 370 121 404 497
rect 628 121 662 497
rect 886 121 920 497
rect 1144 121 1178 497
rect 1402 121 1436 497
rect 1660 121 1694 497
rect 1918 121 1952 497
rect -1952 -435 -1918 -59
rect -1694 -435 -1660 -59
rect -1436 -435 -1402 -59
rect -1178 -435 -1144 -59
rect -920 -435 -886 -59
rect -662 -435 -628 -59
rect -404 -435 -370 -59
rect -146 -435 -112 -59
rect 112 -435 146 -59
rect 370 -435 404 -59
rect 628 -435 662 -59
rect 886 -435 920 -59
rect 1144 -435 1178 -59
rect 1402 -435 1436 -59
rect 1660 -435 1694 -59
rect 1918 -435 1952 -59
<< psubdiff >>
rect -2066 587 -1970 621
rect 1970 587 2066 621
rect -2066 525 -2032 587
rect 2032 525 2066 587
rect -2066 -587 -2032 -525
rect 2032 -587 2066 -525
rect -2066 -621 2066 -587
<< psubdiffcont >>
rect -1970 587 1970 621
rect -2066 -525 -2032 525
rect 2032 -525 2066 525
<< poly >>
rect -1906 509 -1706 535
rect -1648 509 -1448 535
rect -1390 509 -1190 535
rect -1132 509 -932 535
rect -874 509 -674 535
rect -616 509 -416 535
rect -358 509 -158 535
rect -100 509 100 535
rect 158 509 358 535
rect 416 509 616 535
rect 674 509 874 535
rect 932 509 1132 535
rect 1190 509 1390 535
rect 1448 509 1648 535
rect 1706 509 1906 535
rect -1906 71 -1706 109
rect -1906 37 -1890 71
rect -1722 37 -1706 71
rect -1906 21 -1706 37
rect -1648 71 -1448 109
rect -1648 37 -1632 71
rect -1464 37 -1448 71
rect -1648 21 -1448 37
rect -1390 71 -1190 109
rect -1390 37 -1374 71
rect -1206 37 -1190 71
rect -1390 21 -1190 37
rect -1132 71 -932 109
rect -1132 37 -1116 71
rect -948 37 -932 71
rect -1132 21 -932 37
rect -874 71 -674 109
rect -874 37 -858 71
rect -690 37 -674 71
rect -874 21 -674 37
rect -616 71 -416 109
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 109
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 109
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 109
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect 674 71 874 109
rect 674 37 690 71
rect 858 37 874 71
rect 674 21 874 37
rect 932 71 1132 109
rect 932 37 948 71
rect 1116 37 1132 71
rect 932 21 1132 37
rect 1190 71 1390 109
rect 1190 37 1206 71
rect 1374 37 1390 71
rect 1190 21 1390 37
rect 1448 71 1648 109
rect 1448 37 1464 71
rect 1632 37 1648 71
rect 1448 21 1648 37
rect 1706 71 1906 109
rect 1706 37 1722 71
rect 1890 37 1906 71
rect 1706 21 1906 37
rect -1906 -47 -1706 -21
rect -1648 -47 -1448 -21
rect -1390 -47 -1190 -21
rect -1132 -47 -932 -21
rect -874 -47 -674 -21
rect -616 -47 -416 -21
rect -358 -47 -158 -21
rect -100 -47 100 -21
rect 158 -47 358 -21
rect 416 -47 616 -21
rect 674 -47 874 -21
rect 932 -47 1132 -21
rect 1190 -47 1390 -21
rect 1448 -47 1648 -21
rect 1706 -47 1906 -21
rect -1906 -485 -1706 -447
rect -1906 -519 -1890 -485
rect -1722 -519 -1706 -485
rect -1906 -535 -1706 -519
rect -1648 -485 -1448 -447
rect -1648 -519 -1632 -485
rect -1464 -519 -1448 -485
rect -1648 -535 -1448 -519
rect -1390 -485 -1190 -447
rect -1390 -519 -1374 -485
rect -1206 -519 -1190 -485
rect -1390 -535 -1190 -519
rect -1132 -485 -932 -447
rect -1132 -519 -1116 -485
rect -948 -519 -932 -485
rect -1132 -535 -932 -519
rect -874 -485 -674 -447
rect -874 -519 -858 -485
rect -690 -519 -674 -485
rect -874 -535 -674 -519
rect -616 -485 -416 -447
rect -616 -519 -600 -485
rect -432 -519 -416 -485
rect -616 -535 -416 -519
rect -358 -485 -158 -447
rect -358 -519 -342 -485
rect -174 -519 -158 -485
rect -358 -535 -158 -519
rect -100 -485 100 -447
rect -100 -519 -84 -485
rect 84 -519 100 -485
rect -100 -535 100 -519
rect 158 -485 358 -447
rect 158 -519 174 -485
rect 342 -519 358 -485
rect 158 -535 358 -519
rect 416 -485 616 -447
rect 416 -519 432 -485
rect 600 -519 616 -485
rect 416 -535 616 -519
rect 674 -485 874 -447
rect 674 -519 690 -485
rect 858 -519 874 -485
rect 674 -535 874 -519
rect 932 -485 1132 -447
rect 932 -519 948 -485
rect 1116 -519 1132 -485
rect 932 -535 1132 -519
rect 1190 -485 1390 -447
rect 1190 -519 1206 -485
rect 1374 -519 1390 -485
rect 1190 -535 1390 -519
rect 1448 -485 1648 -447
rect 1448 -519 1464 -485
rect 1632 -519 1648 -485
rect 1448 -535 1648 -519
rect 1706 -485 1906 -447
rect 1706 -519 1722 -485
rect 1890 -519 1906 -485
rect 1706 -535 1906 -519
<< polycont >>
rect -1890 37 -1722 71
rect -1632 37 -1464 71
rect -1374 37 -1206 71
rect -1116 37 -948 71
rect -858 37 -690 71
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect 690 37 858 71
rect 948 37 1116 71
rect 1206 37 1374 71
rect 1464 37 1632 71
rect 1722 37 1890 71
rect -1890 -519 -1722 -485
rect -1632 -519 -1464 -485
rect -1374 -519 -1206 -485
rect -1116 -519 -948 -485
rect -858 -519 -690 -485
rect -600 -519 -432 -485
rect -342 -519 -174 -485
rect -84 -519 84 -485
rect 174 -519 342 -485
rect 432 -519 600 -485
rect 690 -519 858 -485
rect 948 -519 1116 -485
rect 1206 -519 1374 -485
rect 1464 -519 1632 -485
rect 1722 -519 1890 -485
<< locali >>
rect -2066 525 -2032 621
rect 2032 525 2066 621
rect -1952 497 -1918 513
rect -1952 105 -1918 121
rect -1694 497 -1660 513
rect -1694 105 -1660 121
rect -1436 497 -1402 513
rect -1436 105 -1402 121
rect -1178 497 -1144 513
rect -1178 105 -1144 121
rect -920 497 -886 513
rect -920 105 -886 121
rect -662 497 -628 513
rect -662 105 -628 121
rect -404 497 -370 513
rect -404 105 -370 121
rect -146 497 -112 513
rect -146 105 -112 121
rect 112 497 146 513
rect 112 105 146 121
rect 370 497 404 513
rect 370 105 404 121
rect 628 497 662 513
rect 628 105 662 121
rect 886 497 920 513
rect 886 105 920 121
rect 1144 497 1178 513
rect 1144 105 1178 121
rect 1402 497 1436 513
rect 1402 105 1436 121
rect 1660 497 1694 513
rect 1660 105 1694 121
rect 1918 497 1952 513
rect 1918 105 1952 121
rect -1906 37 -1890 71
rect -1722 37 -1706 71
rect -1648 37 -1632 71
rect -1464 37 -1448 71
rect -1390 37 -1374 71
rect -1206 37 -1190 71
rect -1132 37 -1116 71
rect -948 37 -932 71
rect -874 37 -858 71
rect -690 37 -674 71
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect 674 37 690 71
rect 858 37 874 71
rect 932 37 948 71
rect 1116 37 1132 71
rect 1190 37 1206 71
rect 1374 37 1390 71
rect 1448 37 1464 71
rect 1632 37 1648 71
rect 1706 37 1722 71
rect 1890 37 1906 71
rect -1952 -59 -1918 -43
rect -1952 -451 -1918 -435
rect -1694 -59 -1660 -43
rect -1694 -451 -1660 -435
rect -1436 -59 -1402 -43
rect -1436 -451 -1402 -435
rect -1178 -59 -1144 -43
rect -1178 -451 -1144 -435
rect -920 -59 -886 -43
rect -920 -451 -886 -435
rect -662 -59 -628 -43
rect -662 -451 -628 -435
rect -404 -59 -370 -43
rect -404 -451 -370 -435
rect -146 -59 -112 -43
rect -146 -451 -112 -435
rect 112 -59 146 -43
rect 112 -451 146 -435
rect 370 -59 404 -43
rect 370 -451 404 -435
rect 628 -59 662 -43
rect 628 -451 662 -435
rect 886 -59 920 -43
rect 886 -451 920 -435
rect 1144 -59 1178 -43
rect 1144 -451 1178 -435
rect 1402 -59 1436 -43
rect 1402 -451 1436 -435
rect 1660 -59 1694 -43
rect 1660 -451 1694 -435
rect 1918 -59 1952 -43
rect 1918 -451 1952 -435
rect -1906 -519 -1890 -485
rect -1722 -519 -1706 -485
rect -1648 -519 -1632 -485
rect -1464 -519 -1448 -485
rect -1390 -519 -1374 -485
rect -1206 -519 -1190 -485
rect -1132 -519 -1116 -485
rect -948 -519 -932 -485
rect -874 -519 -858 -485
rect -690 -519 -674 -485
rect -616 -519 -600 -485
rect -432 -519 -416 -485
rect -358 -519 -342 -485
rect -174 -519 -158 -485
rect -100 -519 -84 -485
rect 84 -519 100 -485
rect 158 -519 174 -485
rect 342 -519 358 -485
rect 416 -519 432 -485
rect 600 -519 616 -485
rect 674 -519 690 -485
rect 858 -519 874 -485
rect 932 -519 948 -485
rect 1116 -519 1132 -485
rect 1190 -519 1206 -485
rect 1374 -519 1390 -485
rect 1448 -519 1464 -485
rect 1632 -519 1648 -485
rect 1706 -519 1722 -485
rect 1890 -519 1906 -485
rect -2066 -621 2066 -587
<< viali >>
rect -2032 587 -1970 621
rect -1970 587 1970 621
rect 1970 587 2032 621
rect -1952 330 -1918 480
rect -1694 138 -1660 288
rect -1436 330 -1402 480
rect -1178 138 -1144 288
rect -920 330 -886 480
rect -662 138 -628 288
rect -404 330 -370 480
rect -146 138 -112 288
rect 112 330 146 480
rect 370 138 404 288
rect 628 330 662 480
rect 886 138 920 288
rect 1144 330 1178 480
rect 1402 138 1436 288
rect 1660 330 1694 480
rect 1918 138 1952 288
rect -1890 37 -1722 71
rect -1632 37 -1464 71
rect -1374 37 -1206 71
rect -1116 37 -948 71
rect -858 37 -690 71
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect 690 37 858 71
rect 948 37 1116 71
rect 1206 37 1374 71
rect 1464 37 1632 71
rect 1722 37 1890 71
rect -2066 -525 -2032 -117
rect -1952 -226 -1918 -76
rect -1694 -418 -1660 -268
rect -1436 -226 -1402 -76
rect -1178 -418 -1144 -268
rect -920 -226 -886 -76
rect -662 -418 -628 -268
rect -404 -226 -370 -76
rect -146 -418 -112 -268
rect 112 -226 146 -76
rect 370 -418 404 -268
rect 628 -226 662 -76
rect 886 -418 920 -268
rect 1144 -226 1178 -76
rect 1402 -418 1436 -268
rect 1660 -226 1694 -76
rect 1918 -418 1952 -268
rect -1890 -519 -1722 -485
rect -1632 -519 -1464 -485
rect -1374 -519 -1206 -485
rect -1116 -519 -948 -485
rect -858 -519 -690 -485
rect -600 -519 -432 -485
rect -342 -519 -174 -485
rect -84 -519 84 -485
rect 174 -519 342 -485
rect 432 -519 600 -485
rect 690 -519 858 -485
rect 948 -519 1116 -485
rect 1206 -519 1374 -485
rect 1464 -519 1632 -485
rect 1722 -519 1890 -485
rect -2066 -587 -2032 -525
rect 2032 -525 2066 -117
rect 2032 -587 2066 -525
<< metal1 >>
rect -2044 621 2044 627
rect -2044 587 -2032 621
rect 2032 587 2044 621
rect -2044 581 2044 587
rect -1958 480 -1912 492
rect -1958 330 -1952 480
rect -1918 330 -1912 480
rect -1958 318 -1912 330
rect -1442 480 -1396 492
rect -1442 330 -1436 480
rect -1402 330 -1396 480
rect -1442 318 -1396 330
rect -926 480 -880 492
rect -926 330 -920 480
rect -886 330 -880 480
rect -926 318 -880 330
rect -410 480 -364 492
rect -410 330 -404 480
rect -370 330 -364 480
rect -410 318 -364 330
rect 106 480 152 492
rect 106 330 112 480
rect 146 330 152 480
rect 106 318 152 330
rect 622 480 668 492
rect 622 330 628 480
rect 662 330 668 480
rect 622 318 668 330
rect 1138 480 1184 492
rect 1138 330 1144 480
rect 1178 330 1184 480
rect 1138 318 1184 330
rect 1654 480 1700 492
rect 1654 330 1660 480
rect 1694 330 1700 480
rect 1654 318 1700 330
rect -1700 288 -1654 300
rect -1700 138 -1694 288
rect -1660 138 -1654 288
rect -1700 126 -1654 138
rect -1184 288 -1138 300
rect -1184 138 -1178 288
rect -1144 138 -1138 288
rect -1184 126 -1138 138
rect -668 288 -622 300
rect -668 138 -662 288
rect -628 138 -622 288
rect -668 126 -622 138
rect -152 288 -106 300
rect -152 138 -146 288
rect -112 138 -106 288
rect -152 126 -106 138
rect 364 288 410 300
rect 364 138 370 288
rect 404 138 410 288
rect 364 126 410 138
rect 880 288 926 300
rect 880 138 886 288
rect 920 138 926 288
rect 880 126 926 138
rect 1396 288 1442 300
rect 1396 138 1402 288
rect 1436 138 1442 288
rect 1396 126 1442 138
rect 1912 288 1958 300
rect 1912 138 1918 288
rect 1952 138 1958 288
rect 1912 126 1958 138
rect -1902 71 -1710 77
rect -1902 37 -1890 71
rect -1722 37 -1710 71
rect -1902 31 -1710 37
rect -1644 71 -1452 77
rect -1644 37 -1632 71
rect -1464 37 -1452 71
rect -1644 31 -1452 37
rect -1386 71 -1194 77
rect -1386 37 -1374 71
rect -1206 37 -1194 71
rect -1386 31 -1194 37
rect -1128 71 -936 77
rect -1128 37 -1116 71
rect -948 37 -936 71
rect -1128 31 -936 37
rect -870 71 -678 77
rect -870 37 -858 71
rect -690 37 -678 71
rect -870 31 -678 37
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect 678 71 870 77
rect 678 37 690 71
rect 858 37 870 71
rect 678 31 870 37
rect 936 71 1128 77
rect 936 37 948 71
rect 1116 37 1128 71
rect 936 31 1128 37
rect 1194 71 1386 77
rect 1194 37 1206 71
rect 1374 37 1386 71
rect 1194 31 1386 37
rect 1452 71 1644 77
rect 1452 37 1464 71
rect 1632 37 1644 71
rect 1452 31 1644 37
rect 1710 71 1902 77
rect 1710 37 1722 71
rect 1890 37 1902 71
rect 1710 31 1902 37
rect -1958 -76 -1912 -64
rect -2072 -117 -2026 -105
rect -2072 -587 -2066 -117
rect -2032 -587 -2026 -117
rect -1958 -226 -1952 -76
rect -1918 -226 -1912 -76
rect -1958 -238 -1912 -226
rect -1442 -76 -1396 -64
rect -1442 -226 -1436 -76
rect -1402 -226 -1396 -76
rect -1442 -238 -1396 -226
rect -926 -76 -880 -64
rect -926 -226 -920 -76
rect -886 -226 -880 -76
rect -926 -238 -880 -226
rect -410 -76 -364 -64
rect -410 -226 -404 -76
rect -370 -226 -364 -76
rect -410 -238 -364 -226
rect 106 -76 152 -64
rect 106 -226 112 -76
rect 146 -226 152 -76
rect 106 -238 152 -226
rect 622 -76 668 -64
rect 622 -226 628 -76
rect 662 -226 668 -76
rect 622 -238 668 -226
rect 1138 -76 1184 -64
rect 1138 -226 1144 -76
rect 1178 -226 1184 -76
rect 1138 -238 1184 -226
rect 1654 -76 1700 -64
rect 1654 -226 1660 -76
rect 1694 -226 1700 -76
rect 1654 -238 1700 -226
rect 2026 -117 2072 -105
rect -1700 -268 -1654 -256
rect -1700 -418 -1694 -268
rect -1660 -418 -1654 -268
rect -1700 -430 -1654 -418
rect -1184 -268 -1138 -256
rect -1184 -418 -1178 -268
rect -1144 -418 -1138 -268
rect -1184 -430 -1138 -418
rect -668 -268 -622 -256
rect -668 -418 -662 -268
rect -628 -418 -622 -268
rect -668 -430 -622 -418
rect -152 -268 -106 -256
rect -152 -418 -146 -268
rect -112 -418 -106 -268
rect -152 -430 -106 -418
rect 364 -268 410 -256
rect 364 -418 370 -268
rect 404 -418 410 -268
rect 364 -430 410 -418
rect 880 -268 926 -256
rect 880 -418 886 -268
rect 920 -418 926 -268
rect 880 -430 926 -418
rect 1396 -268 1442 -256
rect 1396 -418 1402 -268
rect 1436 -418 1442 -268
rect 1396 -430 1442 -418
rect 1912 -268 1958 -256
rect 1912 -418 1918 -268
rect 1952 -418 1958 -268
rect 1912 -430 1958 -418
rect -1902 -485 -1710 -479
rect -1902 -519 -1890 -485
rect -1722 -519 -1710 -485
rect -1902 -525 -1710 -519
rect -1644 -485 -1452 -479
rect -1644 -519 -1632 -485
rect -1464 -519 -1452 -485
rect -1644 -525 -1452 -519
rect -1386 -485 -1194 -479
rect -1386 -519 -1374 -485
rect -1206 -519 -1194 -485
rect -1386 -525 -1194 -519
rect -1128 -485 -936 -479
rect -1128 -519 -1116 -485
rect -948 -519 -936 -485
rect -1128 -525 -936 -519
rect -870 -485 -678 -479
rect -870 -519 -858 -485
rect -690 -519 -678 -485
rect -870 -525 -678 -519
rect -612 -485 -420 -479
rect -612 -519 -600 -485
rect -432 -519 -420 -485
rect -612 -525 -420 -519
rect -354 -485 -162 -479
rect -354 -519 -342 -485
rect -174 -519 -162 -485
rect -354 -525 -162 -519
rect -96 -485 96 -479
rect -96 -519 -84 -485
rect 84 -519 96 -485
rect -96 -525 96 -519
rect 162 -485 354 -479
rect 162 -519 174 -485
rect 342 -519 354 -485
rect 162 -525 354 -519
rect 420 -485 612 -479
rect 420 -519 432 -485
rect 600 -519 612 -485
rect 420 -525 612 -519
rect 678 -485 870 -479
rect 678 -519 690 -485
rect 858 -519 870 -485
rect 678 -525 870 -519
rect 936 -485 1128 -479
rect 936 -519 948 -485
rect 1116 -519 1128 -485
rect 936 -525 1128 -519
rect 1194 -485 1386 -479
rect 1194 -519 1206 -485
rect 1374 -519 1386 -485
rect 1194 -525 1386 -519
rect 1452 -485 1644 -479
rect 1452 -519 1464 -485
rect 1632 -519 1644 -485
rect 1452 -525 1644 -519
rect 1710 -485 1902 -479
rect 1710 -519 1722 -485
rect 1890 -519 1902 -485
rect 1710 -525 1902 -519
rect -2072 -599 -2026 -587
rect 2026 -587 2032 -117
rect 2066 -587 2072 -117
rect 2026 -599 2072 -587
<< properties >>
string FIXED_BBOX -2049 -604 2049 604
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
