magic
tech sky130A
timestamp 1713067979
<< pwell >>
rect -341 -505 341 505
<< nmos >>
rect -243 -400 -143 400
rect -114 -400 -14 400
rect 14 -400 114 400
rect 143 -400 243 400
<< ndiff >>
rect -272 394 -243 400
rect -272 -394 -266 394
rect -249 -394 -243 394
rect -272 -400 -243 -394
rect -143 394 -114 400
rect -143 -394 -137 394
rect -120 -394 -114 394
rect -143 -400 -114 -394
rect -14 394 14 400
rect -14 -394 -8 394
rect 8 -394 14 394
rect -14 -400 14 -394
rect 114 394 143 400
rect 114 -394 120 394
rect 137 -394 143 394
rect 114 -400 143 -394
rect 243 394 272 400
rect 243 -394 249 394
rect 266 -394 272 394
rect 243 -400 272 -394
<< ndiffc >>
rect -266 -394 -249 394
rect -137 -394 -120 394
rect -8 -394 8 394
rect 120 -394 137 394
rect 249 -394 266 394
<< psubdiff >>
rect -323 470 323 487
rect -323 439 -306 470
rect 306 439 323 470
rect -323 -470 -306 -439
rect 306 -470 323 -439
rect -323 -487 -275 -470
rect 275 -487 323 -470
<< psubdiffcont >>
rect -323 -439 -306 439
rect 306 -439 323 439
rect -275 -487 275 -470
<< poly >>
rect -243 436 -143 444
rect -243 419 -235 436
rect -151 419 -143 436
rect -243 400 -143 419
rect -114 436 -14 444
rect -114 419 -106 436
rect -22 419 -14 436
rect -114 400 -14 419
rect 14 436 114 444
rect 14 419 22 436
rect 106 419 114 436
rect 14 400 114 419
rect 143 436 243 444
rect 143 419 151 436
rect 235 419 243 436
rect 143 400 243 419
rect -243 -419 -143 -400
rect -243 -436 -235 -419
rect -151 -436 -143 -419
rect -243 -444 -143 -436
rect -114 -419 -14 -400
rect -114 -436 -106 -419
rect -22 -436 -14 -419
rect -114 -444 -14 -436
rect 14 -419 114 -400
rect 14 -436 22 -419
rect 106 -436 114 -419
rect 14 -444 114 -436
rect 143 -419 243 -400
rect 143 -436 151 -419
rect 235 -436 243 -419
rect 143 -444 243 -436
<< polycont >>
rect -235 419 -151 436
rect -106 419 -22 436
rect 22 419 106 436
rect 151 419 235 436
rect -235 -436 -151 -419
rect -106 -436 -22 -419
rect 22 -436 106 -419
rect 151 -436 235 -419
<< locali >>
rect -323 439 -306 487
rect 306 439 323 487
rect -243 419 -235 436
rect -151 419 -143 436
rect -114 419 -106 436
rect -22 419 -14 436
rect 14 419 22 436
rect 106 419 114 436
rect 143 419 151 436
rect 235 419 243 436
rect -266 394 -249 402
rect -266 -402 -249 -394
rect -137 394 -120 402
rect -137 -402 -120 -394
rect -8 394 8 402
rect -8 -402 8 -394
rect 120 394 137 402
rect 120 -402 137 -394
rect 249 394 266 402
rect 249 -402 266 -394
rect -243 -436 -235 -419
rect -151 -436 -143 -419
rect -114 -436 -106 -419
rect -22 -436 -14 -419
rect 14 -436 22 -419
rect 106 -436 114 -419
rect 143 -436 151 -419
rect 235 -436 243 -419
rect -323 -487 -275 -470
rect 275 -487 323 -470
<< viali >>
rect -306 470 306 487
rect -235 419 -151 436
rect -106 419 -22 436
rect 22 419 106 436
rect 151 419 235 436
rect -323 -439 -306 -94
rect -266 70 -249 385
rect -137 -385 -120 -70
rect -8 70 8 385
rect 120 -385 137 -70
rect 249 70 266 385
rect -235 -436 -151 -419
rect -106 -436 -22 -419
rect 22 -436 106 -419
rect 151 -436 235 -419
rect -323 -470 -306 -439
rect 306 -439 323 -94
rect 306 -470 323 -439
<< metal1 >>
rect -312 487 312 490
rect -312 470 -306 487
rect 306 470 312 487
rect -312 467 312 470
rect -241 436 -145 439
rect -241 419 -235 436
rect -151 419 -145 436
rect -241 416 -145 419
rect -112 436 -16 439
rect -112 419 -106 436
rect -22 419 -16 436
rect -112 416 -16 419
rect 16 436 112 439
rect 16 419 22 436
rect 106 419 112 436
rect 16 416 112 419
rect 145 436 241 439
rect 145 419 151 436
rect 235 419 241 436
rect 145 416 241 419
rect -269 385 -246 391
rect -269 70 -266 385
rect -249 70 -246 385
rect -269 64 -246 70
rect -11 385 11 391
rect -11 70 -8 385
rect 8 70 11 385
rect -11 64 11 70
rect 246 385 269 391
rect 246 70 249 385
rect 266 70 269 385
rect 246 64 269 70
rect -140 -70 -117 -64
rect -326 -94 -303 -88
rect -326 -470 -323 -94
rect -306 -470 -303 -94
rect -140 -385 -137 -70
rect -120 -385 -117 -70
rect -140 -391 -117 -385
rect 117 -70 140 -64
rect 117 -385 120 -70
rect 137 -385 140 -70
rect 117 -391 140 -385
rect 303 -94 326 -88
rect -241 -419 -145 -416
rect -241 -436 -235 -419
rect -151 -436 -145 -419
rect -241 -439 -145 -436
rect -112 -419 -16 -416
rect -112 -436 -106 -419
rect -22 -436 -16 -419
rect -112 -439 -16 -436
rect 16 -419 112 -416
rect 16 -436 22 -419
rect 106 -436 112 -419
rect 16 -439 112 -436
rect 145 -419 241 -416
rect 145 -436 151 -419
rect 235 -436 241 -419
rect 145 -439 241 -436
rect -326 -476 -303 -470
rect 303 -470 306 -94
rect 323 -470 326 -94
rect 303 -476 326 -470
<< properties >>
string FIXED_BBOX -315 -478 315 478
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr +40 viagl +40 viagt 100
<< end >>
