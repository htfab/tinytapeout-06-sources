magic
tech sky130A
timestamp 1713539272
<< pwell >>
rect -148 -905 148 905
<< nmoslvt >>
rect -50 -800 50 800
<< ndiff >>
rect -79 794 -50 800
rect -79 -794 -73 794
rect -56 -794 -50 794
rect -79 -800 -50 -794
rect 50 794 79 800
rect 50 -794 56 794
rect 73 -794 79 794
rect 50 -800 79 -794
<< ndiffc >>
rect -73 -794 -56 794
rect 56 -794 73 794
<< psubdiff >>
rect -130 870 -82 887
rect 82 870 130 887
rect -130 839 -113 870
rect 113 839 130 870
rect -130 -870 -113 -839
rect 113 -870 130 -839
rect -130 -887 -82 -870
rect 82 -887 130 -870
<< psubdiffcont >>
rect -82 870 82 887
rect -130 -839 -113 839
rect 113 -839 130 839
rect -82 -887 82 -870
<< poly >>
rect -50 836 50 844
rect -50 819 -42 836
rect 42 819 50 836
rect -50 800 50 819
rect -50 -819 50 -800
rect -50 -836 -42 -819
rect 42 -836 50 -819
rect -50 -844 50 -836
<< polycont >>
rect -42 819 42 836
rect -42 -836 42 -819
<< locali >>
rect -130 870 -82 887
rect 82 870 130 887
rect -130 839 -113 870
rect 113 839 130 870
rect -50 819 -42 836
rect 42 819 50 836
rect -73 794 -56 802
rect -73 -802 -56 -794
rect 56 794 73 802
rect 56 -802 73 -794
rect -50 -836 -42 -819
rect 42 -836 50 -819
rect -130 -870 -113 -839
rect 113 -870 130 -839
rect -130 -887 -82 -870
rect 82 -887 130 -870
<< viali >>
rect -42 819 42 836
rect -73 -794 -56 794
rect 56 -794 73 794
rect -42 -836 42 -819
<< metal1 >>
rect -48 836 48 839
rect -48 819 -42 836
rect 42 819 48 836
rect -48 816 48 819
rect -76 794 -53 800
rect -76 -794 -73 794
rect -56 -794 -53 794
rect -76 -800 -53 -794
rect 53 794 76 800
rect 53 -794 56 794
rect 73 -794 76 794
rect 53 -800 76 -794
rect -48 -819 48 -816
rect -48 -836 -42 -819
rect 42 -836 48 -819
rect -48 -839 48 -836
<< properties >>
string FIXED_BBOX -121 -878 121 878
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 16.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
