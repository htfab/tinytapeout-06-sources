** sch_path: /home/dsatizabal/tt06-fet-opamp/xschem/opamp.sch
.subckt opamp VDD ZREF vin_n vin_p Vout VGND
*.PININFO vin_n:I vin_p:I Vout:O VDD:B ZREF:B VGND:B
XM1 net1 vin_n net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM2 net2 vin_p net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM3 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 m=1
XM4 net2 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 m=1
XM5 net3 VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM7 Vout VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM8 ZREF VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM9 net4 VDD net2 VGND sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 m=1
XC1 net4 Vout sky130_fd_pr__cap_mim_m3_1 W=17.55 L=15 m=1
XM6 Vout net2 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 m=1
XR1 ZREF VDD VGND sky130_fd_pr__res_generic_nd W=1 L=5 mult=1 m=1
XR2 VGND ZREF VGND sky130_fd_pr__res_generic_nd W=1 L=5 mult=1 m=1
.ends
.end
