magic
tech sky130A
magscale 1 2
timestamp 1713448216
<< nwell >>
rect -296 -16871 296 16871
<< pmos >>
rect -100 14652 100 16652
rect -100 12416 100 14416
rect -100 10180 100 12180
rect -100 7944 100 9944
rect -100 5708 100 7708
rect -100 3472 100 5472
rect -100 1236 100 3236
rect -100 -1000 100 1000
rect -100 -3236 100 -1236
rect -100 -5472 100 -3472
rect -100 -7708 100 -5708
rect -100 -9944 100 -7944
rect -100 -12180 100 -10180
rect -100 -14416 100 -12416
rect -100 -16652 100 -14652
<< pdiff >>
rect -158 16640 -100 16652
rect -158 14664 -146 16640
rect -112 14664 -100 16640
rect -158 14652 -100 14664
rect 100 16640 158 16652
rect 100 14664 112 16640
rect 146 14664 158 16640
rect 100 14652 158 14664
rect -158 14404 -100 14416
rect -158 12428 -146 14404
rect -112 12428 -100 14404
rect -158 12416 -100 12428
rect 100 14404 158 14416
rect 100 12428 112 14404
rect 146 12428 158 14404
rect 100 12416 158 12428
rect -158 12168 -100 12180
rect -158 10192 -146 12168
rect -112 10192 -100 12168
rect -158 10180 -100 10192
rect 100 12168 158 12180
rect 100 10192 112 12168
rect 146 10192 158 12168
rect 100 10180 158 10192
rect -158 9932 -100 9944
rect -158 7956 -146 9932
rect -112 7956 -100 9932
rect -158 7944 -100 7956
rect 100 9932 158 9944
rect 100 7956 112 9932
rect 146 7956 158 9932
rect 100 7944 158 7956
rect -158 7696 -100 7708
rect -158 5720 -146 7696
rect -112 5720 -100 7696
rect -158 5708 -100 5720
rect 100 7696 158 7708
rect 100 5720 112 7696
rect 146 5720 158 7696
rect 100 5708 158 5720
rect -158 5460 -100 5472
rect -158 3484 -146 5460
rect -112 3484 -100 5460
rect -158 3472 -100 3484
rect 100 5460 158 5472
rect 100 3484 112 5460
rect 146 3484 158 5460
rect 100 3472 158 3484
rect -158 3224 -100 3236
rect -158 1248 -146 3224
rect -112 1248 -100 3224
rect -158 1236 -100 1248
rect 100 3224 158 3236
rect 100 1248 112 3224
rect 146 1248 158 3224
rect 100 1236 158 1248
rect -158 988 -100 1000
rect -158 -988 -146 988
rect -112 -988 -100 988
rect -158 -1000 -100 -988
rect 100 988 158 1000
rect 100 -988 112 988
rect 146 -988 158 988
rect 100 -1000 158 -988
rect -158 -1248 -100 -1236
rect -158 -3224 -146 -1248
rect -112 -3224 -100 -1248
rect -158 -3236 -100 -3224
rect 100 -1248 158 -1236
rect 100 -3224 112 -1248
rect 146 -3224 158 -1248
rect 100 -3236 158 -3224
rect -158 -3484 -100 -3472
rect -158 -5460 -146 -3484
rect -112 -5460 -100 -3484
rect -158 -5472 -100 -5460
rect 100 -3484 158 -3472
rect 100 -5460 112 -3484
rect 146 -5460 158 -3484
rect 100 -5472 158 -5460
rect -158 -5720 -100 -5708
rect -158 -7696 -146 -5720
rect -112 -7696 -100 -5720
rect -158 -7708 -100 -7696
rect 100 -5720 158 -5708
rect 100 -7696 112 -5720
rect 146 -7696 158 -5720
rect 100 -7708 158 -7696
rect -158 -7956 -100 -7944
rect -158 -9932 -146 -7956
rect -112 -9932 -100 -7956
rect -158 -9944 -100 -9932
rect 100 -7956 158 -7944
rect 100 -9932 112 -7956
rect 146 -9932 158 -7956
rect 100 -9944 158 -9932
rect -158 -10192 -100 -10180
rect -158 -12168 -146 -10192
rect -112 -12168 -100 -10192
rect -158 -12180 -100 -12168
rect 100 -10192 158 -10180
rect 100 -12168 112 -10192
rect 146 -12168 158 -10192
rect 100 -12180 158 -12168
rect -158 -12428 -100 -12416
rect -158 -14404 -146 -12428
rect -112 -14404 -100 -12428
rect -158 -14416 -100 -14404
rect 100 -12428 158 -12416
rect 100 -14404 112 -12428
rect 146 -14404 158 -12428
rect 100 -14416 158 -14404
rect -158 -14664 -100 -14652
rect -158 -16640 -146 -14664
rect -112 -16640 -100 -14664
rect -158 -16652 -100 -16640
rect 100 -14664 158 -14652
rect 100 -16640 112 -14664
rect 146 -16640 158 -14664
rect 100 -16652 158 -16640
<< pdiffc >>
rect -146 14664 -112 16640
rect 112 14664 146 16640
rect -146 12428 -112 14404
rect 112 12428 146 14404
rect -146 10192 -112 12168
rect 112 10192 146 12168
rect -146 7956 -112 9932
rect 112 7956 146 9932
rect -146 5720 -112 7696
rect 112 5720 146 7696
rect -146 3484 -112 5460
rect 112 3484 146 5460
rect -146 1248 -112 3224
rect 112 1248 146 3224
rect -146 -988 -112 988
rect 112 -988 146 988
rect -146 -3224 -112 -1248
rect 112 -3224 146 -1248
rect -146 -5460 -112 -3484
rect 112 -5460 146 -3484
rect -146 -7696 -112 -5720
rect 112 -7696 146 -5720
rect -146 -9932 -112 -7956
rect 112 -9932 146 -7956
rect -146 -12168 -112 -10192
rect 112 -12168 146 -10192
rect -146 -14404 -112 -12428
rect 112 -14404 146 -12428
rect -146 -16640 -112 -14664
rect 112 -16640 146 -14664
<< nsubdiff >>
rect -260 16801 -164 16835
rect 164 16801 260 16835
rect -260 16739 -226 16801
rect 226 16739 260 16801
rect -260 -16801 -226 -16739
rect 226 -16801 260 -16739
rect -260 -16835 -164 -16801
rect 164 -16835 260 -16801
<< nsubdiffcont >>
rect -164 16801 164 16835
rect -260 -16739 -226 16739
rect 226 -16739 260 16739
rect -164 -16835 164 -16801
<< poly >>
rect -100 16733 100 16749
rect -100 16699 -84 16733
rect 84 16699 100 16733
rect -100 16652 100 16699
rect -100 14605 100 14652
rect -100 14571 -84 14605
rect 84 14571 100 14605
rect -100 14555 100 14571
rect -100 14497 100 14513
rect -100 14463 -84 14497
rect 84 14463 100 14497
rect -100 14416 100 14463
rect -100 12369 100 12416
rect -100 12335 -84 12369
rect 84 12335 100 12369
rect -100 12319 100 12335
rect -100 12261 100 12277
rect -100 12227 -84 12261
rect 84 12227 100 12261
rect -100 12180 100 12227
rect -100 10133 100 10180
rect -100 10099 -84 10133
rect 84 10099 100 10133
rect -100 10083 100 10099
rect -100 10025 100 10041
rect -100 9991 -84 10025
rect 84 9991 100 10025
rect -100 9944 100 9991
rect -100 7897 100 7944
rect -100 7863 -84 7897
rect 84 7863 100 7897
rect -100 7847 100 7863
rect -100 7789 100 7805
rect -100 7755 -84 7789
rect 84 7755 100 7789
rect -100 7708 100 7755
rect -100 5661 100 5708
rect -100 5627 -84 5661
rect 84 5627 100 5661
rect -100 5611 100 5627
rect -100 5553 100 5569
rect -100 5519 -84 5553
rect 84 5519 100 5553
rect -100 5472 100 5519
rect -100 3425 100 3472
rect -100 3391 -84 3425
rect 84 3391 100 3425
rect -100 3375 100 3391
rect -100 3317 100 3333
rect -100 3283 -84 3317
rect 84 3283 100 3317
rect -100 3236 100 3283
rect -100 1189 100 1236
rect -100 1155 -84 1189
rect 84 1155 100 1189
rect -100 1139 100 1155
rect -100 1081 100 1097
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -100 1000 100 1047
rect -100 -1047 100 -1000
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1097 100 -1081
rect -100 -1155 100 -1139
rect -100 -1189 -84 -1155
rect 84 -1189 100 -1155
rect -100 -1236 100 -1189
rect -100 -3283 100 -3236
rect -100 -3317 -84 -3283
rect 84 -3317 100 -3283
rect -100 -3333 100 -3317
rect -100 -3391 100 -3375
rect -100 -3425 -84 -3391
rect 84 -3425 100 -3391
rect -100 -3472 100 -3425
rect -100 -5519 100 -5472
rect -100 -5553 -84 -5519
rect 84 -5553 100 -5519
rect -100 -5569 100 -5553
rect -100 -5627 100 -5611
rect -100 -5661 -84 -5627
rect 84 -5661 100 -5627
rect -100 -5708 100 -5661
rect -100 -7755 100 -7708
rect -100 -7789 -84 -7755
rect 84 -7789 100 -7755
rect -100 -7805 100 -7789
rect -100 -7863 100 -7847
rect -100 -7897 -84 -7863
rect 84 -7897 100 -7863
rect -100 -7944 100 -7897
rect -100 -9991 100 -9944
rect -100 -10025 -84 -9991
rect 84 -10025 100 -9991
rect -100 -10041 100 -10025
rect -100 -10099 100 -10083
rect -100 -10133 -84 -10099
rect 84 -10133 100 -10099
rect -100 -10180 100 -10133
rect -100 -12227 100 -12180
rect -100 -12261 -84 -12227
rect 84 -12261 100 -12227
rect -100 -12277 100 -12261
rect -100 -12335 100 -12319
rect -100 -12369 -84 -12335
rect 84 -12369 100 -12335
rect -100 -12416 100 -12369
rect -100 -14463 100 -14416
rect -100 -14497 -84 -14463
rect 84 -14497 100 -14463
rect -100 -14513 100 -14497
rect -100 -14571 100 -14555
rect -100 -14605 -84 -14571
rect 84 -14605 100 -14571
rect -100 -14652 100 -14605
rect -100 -16699 100 -16652
rect -100 -16733 -84 -16699
rect 84 -16733 100 -16699
rect -100 -16749 100 -16733
<< polycont >>
rect -84 16699 84 16733
rect -84 14571 84 14605
rect -84 14463 84 14497
rect -84 12335 84 12369
rect -84 12227 84 12261
rect -84 10099 84 10133
rect -84 9991 84 10025
rect -84 7863 84 7897
rect -84 7755 84 7789
rect -84 5627 84 5661
rect -84 5519 84 5553
rect -84 3391 84 3425
rect -84 3283 84 3317
rect -84 1155 84 1189
rect -84 1047 84 1081
rect -84 -1081 84 -1047
rect -84 -1189 84 -1155
rect -84 -3317 84 -3283
rect -84 -3425 84 -3391
rect -84 -5553 84 -5519
rect -84 -5661 84 -5627
rect -84 -7789 84 -7755
rect -84 -7897 84 -7863
rect -84 -10025 84 -9991
rect -84 -10133 84 -10099
rect -84 -12261 84 -12227
rect -84 -12369 84 -12335
rect -84 -14497 84 -14463
rect -84 -14605 84 -14571
rect -84 -16733 84 -16699
<< locali >>
rect -260 16801 -164 16835
rect 164 16801 260 16835
rect -260 16739 -226 16801
rect 226 16739 260 16801
rect -100 16699 -84 16733
rect 84 16699 100 16733
rect -146 16640 -112 16656
rect -146 14648 -112 14664
rect 112 16640 146 16656
rect 112 14648 146 14664
rect -100 14571 -84 14605
rect 84 14571 100 14605
rect -100 14463 -84 14497
rect 84 14463 100 14497
rect -146 14404 -112 14420
rect -146 12412 -112 12428
rect 112 14404 146 14420
rect 112 12412 146 12428
rect -100 12335 -84 12369
rect 84 12335 100 12369
rect -100 12227 -84 12261
rect 84 12227 100 12261
rect -146 12168 -112 12184
rect -146 10176 -112 10192
rect 112 12168 146 12184
rect 112 10176 146 10192
rect -100 10099 -84 10133
rect 84 10099 100 10133
rect -100 9991 -84 10025
rect 84 9991 100 10025
rect -146 9932 -112 9948
rect -146 7940 -112 7956
rect 112 9932 146 9948
rect 112 7940 146 7956
rect -100 7863 -84 7897
rect 84 7863 100 7897
rect -100 7755 -84 7789
rect 84 7755 100 7789
rect -146 7696 -112 7712
rect -146 5704 -112 5720
rect 112 7696 146 7712
rect 112 5704 146 5720
rect -100 5627 -84 5661
rect 84 5627 100 5661
rect -100 5519 -84 5553
rect 84 5519 100 5553
rect -146 5460 -112 5476
rect -146 3468 -112 3484
rect 112 5460 146 5476
rect 112 3468 146 3484
rect -100 3391 -84 3425
rect 84 3391 100 3425
rect -100 3283 -84 3317
rect 84 3283 100 3317
rect -146 3224 -112 3240
rect -146 1232 -112 1248
rect 112 3224 146 3240
rect 112 1232 146 1248
rect -100 1155 -84 1189
rect 84 1155 100 1189
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -146 988 -112 1004
rect -146 -1004 -112 -988
rect 112 988 146 1004
rect 112 -1004 146 -988
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1189 -84 -1155
rect 84 -1189 100 -1155
rect -146 -1248 -112 -1232
rect -146 -3240 -112 -3224
rect 112 -1248 146 -1232
rect 112 -3240 146 -3224
rect -100 -3317 -84 -3283
rect 84 -3317 100 -3283
rect -100 -3425 -84 -3391
rect 84 -3425 100 -3391
rect -146 -3484 -112 -3468
rect -146 -5476 -112 -5460
rect 112 -3484 146 -3468
rect 112 -5476 146 -5460
rect -100 -5553 -84 -5519
rect 84 -5553 100 -5519
rect -100 -5661 -84 -5627
rect 84 -5661 100 -5627
rect -146 -5720 -112 -5704
rect -146 -7712 -112 -7696
rect 112 -5720 146 -5704
rect 112 -7712 146 -7696
rect -100 -7789 -84 -7755
rect 84 -7789 100 -7755
rect -100 -7897 -84 -7863
rect 84 -7897 100 -7863
rect -146 -7956 -112 -7940
rect -146 -9948 -112 -9932
rect 112 -7956 146 -7940
rect 112 -9948 146 -9932
rect -100 -10025 -84 -9991
rect 84 -10025 100 -9991
rect -100 -10133 -84 -10099
rect 84 -10133 100 -10099
rect -146 -10192 -112 -10176
rect -146 -12184 -112 -12168
rect 112 -10192 146 -10176
rect 112 -12184 146 -12168
rect -100 -12261 -84 -12227
rect 84 -12261 100 -12227
rect -100 -12369 -84 -12335
rect 84 -12369 100 -12335
rect -146 -12428 -112 -12412
rect -146 -14420 -112 -14404
rect 112 -12428 146 -12412
rect 112 -14420 146 -14404
rect -100 -14497 -84 -14463
rect 84 -14497 100 -14463
rect -100 -14605 -84 -14571
rect 84 -14605 100 -14571
rect -146 -14664 -112 -14648
rect -146 -16656 -112 -16640
rect 112 -14664 146 -14648
rect 112 -16656 146 -16640
rect -100 -16733 -84 -16699
rect 84 -16733 100 -16699
rect -260 -16801 -226 -16739
rect 226 -16801 260 -16739
rect -260 -16835 -164 -16801
rect 164 -16835 260 -16801
<< viali >>
rect -84 16699 84 16733
rect -146 14664 -112 16640
rect 112 14664 146 16640
rect -84 14571 84 14605
rect -84 14463 84 14497
rect -146 12428 -112 14404
rect 112 12428 146 14404
rect -84 12335 84 12369
rect -84 12227 84 12261
rect -146 10192 -112 12168
rect 112 10192 146 12168
rect -84 10099 84 10133
rect -84 9991 84 10025
rect -146 7956 -112 9932
rect 112 7956 146 9932
rect -84 7863 84 7897
rect -84 7755 84 7789
rect -146 5720 -112 7696
rect 112 5720 146 7696
rect -84 5627 84 5661
rect -84 5519 84 5553
rect -146 3484 -112 5460
rect 112 3484 146 5460
rect -84 3391 84 3425
rect -84 3283 84 3317
rect -146 1248 -112 3224
rect 112 1248 146 3224
rect -84 1155 84 1189
rect -84 1047 84 1081
rect -146 -988 -112 988
rect 112 -988 146 988
rect -84 -1081 84 -1047
rect -84 -1189 84 -1155
rect -146 -3224 -112 -1248
rect 112 -3224 146 -1248
rect -84 -3317 84 -3283
rect -84 -3425 84 -3391
rect -146 -5460 -112 -3484
rect 112 -5460 146 -3484
rect -84 -5553 84 -5519
rect -84 -5661 84 -5627
rect -146 -7696 -112 -5720
rect 112 -7696 146 -5720
rect -84 -7789 84 -7755
rect -84 -7897 84 -7863
rect -146 -9932 -112 -7956
rect 112 -9932 146 -7956
rect -84 -10025 84 -9991
rect -84 -10133 84 -10099
rect -146 -12168 -112 -10192
rect 112 -12168 146 -10192
rect -84 -12261 84 -12227
rect -84 -12369 84 -12335
rect -146 -14404 -112 -12428
rect 112 -14404 146 -12428
rect -84 -14497 84 -14463
rect -84 -14605 84 -14571
rect -146 -16640 -112 -14664
rect 112 -16640 146 -14664
rect -84 -16733 84 -16699
<< metal1 >>
rect -96 16733 96 16739
rect -96 16699 -84 16733
rect 84 16699 96 16733
rect -96 16693 96 16699
rect -152 16640 -106 16652
rect -152 14664 -146 16640
rect -112 14664 -106 16640
rect -152 14652 -106 14664
rect 106 16640 152 16652
rect 106 14664 112 16640
rect 146 14664 152 16640
rect 106 14652 152 14664
rect -96 14605 96 14611
rect -96 14571 -84 14605
rect 84 14571 96 14605
rect -96 14565 96 14571
rect -96 14497 96 14503
rect -96 14463 -84 14497
rect 84 14463 96 14497
rect -96 14457 96 14463
rect -152 14404 -106 14416
rect -152 12428 -146 14404
rect -112 12428 -106 14404
rect -152 12416 -106 12428
rect 106 14404 152 14416
rect 106 12428 112 14404
rect 146 12428 152 14404
rect 106 12416 152 12428
rect -96 12369 96 12375
rect -96 12335 -84 12369
rect 84 12335 96 12369
rect -96 12329 96 12335
rect -96 12261 96 12267
rect -96 12227 -84 12261
rect 84 12227 96 12261
rect -96 12221 96 12227
rect -152 12168 -106 12180
rect -152 10192 -146 12168
rect -112 10192 -106 12168
rect -152 10180 -106 10192
rect 106 12168 152 12180
rect 106 10192 112 12168
rect 146 10192 152 12168
rect 106 10180 152 10192
rect -96 10133 96 10139
rect -96 10099 -84 10133
rect 84 10099 96 10133
rect -96 10093 96 10099
rect -96 10025 96 10031
rect -96 9991 -84 10025
rect 84 9991 96 10025
rect -96 9985 96 9991
rect -152 9932 -106 9944
rect -152 7956 -146 9932
rect -112 7956 -106 9932
rect -152 7944 -106 7956
rect 106 9932 152 9944
rect 106 7956 112 9932
rect 146 7956 152 9932
rect 106 7944 152 7956
rect -96 7897 96 7903
rect -96 7863 -84 7897
rect 84 7863 96 7897
rect -96 7857 96 7863
rect -96 7789 96 7795
rect -96 7755 -84 7789
rect 84 7755 96 7789
rect -96 7749 96 7755
rect -152 7696 -106 7708
rect -152 5720 -146 7696
rect -112 5720 -106 7696
rect -152 5708 -106 5720
rect 106 7696 152 7708
rect 106 5720 112 7696
rect 146 5720 152 7696
rect 106 5708 152 5720
rect -96 5661 96 5667
rect -96 5627 -84 5661
rect 84 5627 96 5661
rect -96 5621 96 5627
rect -96 5553 96 5559
rect -96 5519 -84 5553
rect 84 5519 96 5553
rect -96 5513 96 5519
rect -152 5460 -106 5472
rect -152 3484 -146 5460
rect -112 3484 -106 5460
rect -152 3472 -106 3484
rect 106 5460 152 5472
rect 106 3484 112 5460
rect 146 3484 152 5460
rect 106 3472 152 3484
rect -96 3425 96 3431
rect -96 3391 -84 3425
rect 84 3391 96 3425
rect -96 3385 96 3391
rect -96 3317 96 3323
rect -96 3283 -84 3317
rect 84 3283 96 3317
rect -96 3277 96 3283
rect -152 3224 -106 3236
rect -152 1248 -146 3224
rect -112 1248 -106 3224
rect -152 1236 -106 1248
rect 106 3224 152 3236
rect 106 1248 112 3224
rect 146 1248 152 3224
rect 106 1236 152 1248
rect -96 1189 96 1195
rect -96 1155 -84 1189
rect 84 1155 96 1189
rect -96 1149 96 1155
rect -96 1081 96 1087
rect -96 1047 -84 1081
rect 84 1047 96 1081
rect -96 1041 96 1047
rect -152 988 -106 1000
rect -152 -988 -146 988
rect -112 -988 -106 988
rect -152 -1000 -106 -988
rect 106 988 152 1000
rect 106 -988 112 988
rect 146 -988 152 988
rect 106 -1000 152 -988
rect -96 -1047 96 -1041
rect -96 -1081 -84 -1047
rect 84 -1081 96 -1047
rect -96 -1087 96 -1081
rect -96 -1155 96 -1149
rect -96 -1189 -84 -1155
rect 84 -1189 96 -1155
rect -96 -1195 96 -1189
rect -152 -1248 -106 -1236
rect -152 -3224 -146 -1248
rect -112 -3224 -106 -1248
rect -152 -3236 -106 -3224
rect 106 -1248 152 -1236
rect 106 -3224 112 -1248
rect 146 -3224 152 -1248
rect 106 -3236 152 -3224
rect -96 -3283 96 -3277
rect -96 -3317 -84 -3283
rect 84 -3317 96 -3283
rect -96 -3323 96 -3317
rect -96 -3391 96 -3385
rect -96 -3425 -84 -3391
rect 84 -3425 96 -3391
rect -96 -3431 96 -3425
rect -152 -3484 -106 -3472
rect -152 -5460 -146 -3484
rect -112 -5460 -106 -3484
rect -152 -5472 -106 -5460
rect 106 -3484 152 -3472
rect 106 -5460 112 -3484
rect 146 -5460 152 -3484
rect 106 -5472 152 -5460
rect -96 -5519 96 -5513
rect -96 -5553 -84 -5519
rect 84 -5553 96 -5519
rect -96 -5559 96 -5553
rect -96 -5627 96 -5621
rect -96 -5661 -84 -5627
rect 84 -5661 96 -5627
rect -96 -5667 96 -5661
rect -152 -5720 -106 -5708
rect -152 -7696 -146 -5720
rect -112 -7696 -106 -5720
rect -152 -7708 -106 -7696
rect 106 -5720 152 -5708
rect 106 -7696 112 -5720
rect 146 -7696 152 -5720
rect 106 -7708 152 -7696
rect -96 -7755 96 -7749
rect -96 -7789 -84 -7755
rect 84 -7789 96 -7755
rect -96 -7795 96 -7789
rect -96 -7863 96 -7857
rect -96 -7897 -84 -7863
rect 84 -7897 96 -7863
rect -96 -7903 96 -7897
rect -152 -7956 -106 -7944
rect -152 -9932 -146 -7956
rect -112 -9932 -106 -7956
rect -152 -9944 -106 -9932
rect 106 -7956 152 -7944
rect 106 -9932 112 -7956
rect 146 -9932 152 -7956
rect 106 -9944 152 -9932
rect -96 -9991 96 -9985
rect -96 -10025 -84 -9991
rect 84 -10025 96 -9991
rect -96 -10031 96 -10025
rect -96 -10099 96 -10093
rect -96 -10133 -84 -10099
rect 84 -10133 96 -10099
rect -96 -10139 96 -10133
rect -152 -10192 -106 -10180
rect -152 -12168 -146 -10192
rect -112 -12168 -106 -10192
rect -152 -12180 -106 -12168
rect 106 -10192 152 -10180
rect 106 -12168 112 -10192
rect 146 -12168 152 -10192
rect 106 -12180 152 -12168
rect -96 -12227 96 -12221
rect -96 -12261 -84 -12227
rect 84 -12261 96 -12227
rect -96 -12267 96 -12261
rect -96 -12335 96 -12329
rect -96 -12369 -84 -12335
rect 84 -12369 96 -12335
rect -96 -12375 96 -12369
rect -152 -12428 -106 -12416
rect -152 -14404 -146 -12428
rect -112 -14404 -106 -12428
rect -152 -14416 -106 -14404
rect 106 -12428 152 -12416
rect 106 -14404 112 -12428
rect 146 -14404 152 -12428
rect 106 -14416 152 -14404
rect -96 -14463 96 -14457
rect -96 -14497 -84 -14463
rect 84 -14497 96 -14463
rect -96 -14503 96 -14497
rect -96 -14571 96 -14565
rect -96 -14605 -84 -14571
rect 84 -14605 96 -14571
rect -96 -14611 96 -14605
rect -152 -14664 -106 -14652
rect -152 -16640 -146 -14664
rect -112 -16640 -106 -14664
rect -152 -16652 -106 -16640
rect 106 -14664 152 -14652
rect 106 -16640 112 -14664
rect 146 -16640 152 -14664
rect 106 -16652 152 -16640
rect -96 -16699 96 -16693
rect -96 -16733 -84 -16699
rect 84 -16733 96 -16699
rect -96 -16739 96 -16733
<< properties >>
string FIXED_BBOX -243 -16818 243 16818
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 15 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
